BZh91AY&SY�B�	�߀ryg����������`�~    �    m��� (     �  ��{�B�J%	JR�*��8��^�	��K��J�C��^o9�(���s�V;���@��B�wСE !�IT�eƎ�C�Wu� 
us�� |}����E9�s�����T/|w�ύ�4t{f���>���|�. x>���4P�q��cB�c���� :��(��q�r� yh�����Цq� Q����v^4Q�9��N���  /GL�\��W9�(���J U@
P              EH��2�)=S&���44�1����R#*���&�4�a12410jy�$
� 0#&� b`z5RH���       
Q24�i���4�bzL�$yA&�ڢ!)�����x�M��� �;���|�O��}���N�A	?��>�"$�quD T|QD=Ϊ�����n�(#�T1���?�i�~7������8~n�Ӂ�z�M|ߍ�!��=�a��v߯3N࿟���v�}�������?��� *���C�ܱф9�AU@�����UG��S!3*�.������ገ ���
�'=����)�`�׆��٦����U�~����
d�����)��֍
Y�䲯jBi  #�w�p*P���������ߥ3����>�8n��;�;��@7�������_5��yvt�����7wwh-�
¡X((,�wwwv�5
��B�w�X((pq���AB܆�Pnb
�A`��Vq�!X[n���B�V���VۡnB���V

j��V��m�B��(+p-��*
DB�t+PPX(,

����(,x�B���T7qx\���*
���AB����Aa�6ۻB܅B��
"�B�PP���
�A`��
�aP�q�+
��CPXT+8�.�*�wl*

�ATۡm� �XT*q
!Xj
E���q����
�`�P�PPXT8¡XV�b��-�+
�aP�V
��
�����
�aP��-��B��B��V
��P�*�[m�P�*���*
�9Pn��*p*�-��a�!P�+B��T8�*!m�hT
��(,B���ΐ�Ht��((%�T

�j������
�aP�6�aP�q��
�A�*

�m�+
�aPPX(%�m�t I�sd�Ի��+����˩�
�qA����ä:a�!XR�T+�baP����5�b�B܅A�%LL�P�q���T
��B�M������
�8���°�7����m��ۨj�P�*
¡K�^8�B��m��AAaP�[y�
C��T�P�*"��aP�j�XR�[m��B���AT-��+r�����B�PPXT*��1��`�PF�C[��n�
0�[m��ۻ�묇L:���!P�*���P�7-�
�AaP�XT)p��1�B��)p+
��B��
¡XV����aP�%B�
�B��w�C�-����]d�����v�L5
¡P��VP�V
0�T(¡P�\
�¡XT-��
�T*��
�B�D�
�Q
�aP�*
��
�T+
!XQ�B��V׈a����B�XQ�B�B����,-�Tn^`�P�-�T+
��B��VB�XT*m��¡XT*�B�1�T+B��%��*Aj
¡XQ
!XQ
�~������ݰ�T��V
 �
�\��-��ШV
�-��ݡnT+B�F
�^7�`�nB��X(T9�]�2�V
�.B������j
J
Z�%�hh)4�仒��   �.K�B��[��n�������������t���O��OY�:�_��Y;�|y��:?l=���rO�9<�.�/�f|n@w-��6w`s��hs۪g^�h����݄�@A8,���� �&my����FiS��L�Ur���b��/RqŽ;�\�[��!�Z�������q�p:��(�ND�QhX�i�bLC�A�y\��6.TA�xi�q�8�a��a���Lࡈ%# �Ub�!H���s�6mN5<'ė��^��P��;�t�bk ��~J��:��3"&L�\�hG��R�=>��d���7�P�0��OE�5�@��h�=8%��B��s"c��$�R-��"/�ż�SǢ�J_��A8���Xj�'� c���Vn�PS�N������uF���t�"�T�UA�X��U,x�T��H��4�#Bn�74��}���yf�ݥJ�.��I>�(��MML�S����p�"�J��#M�8��Bļ�u�9��(c+#.2br��̡�����Zd���j&���{Ö]H�"&&C�s�nd)�y�up�Fh'jOt��3SJB���C�.�7sx��[��ZyF>n����GԽ�w����j��.g%�1j5FiM`W�N�&2�K���62Մ�O6T]�uss"q�=ӽ,� FL��J^��6mɃC.���B�`�dEVfd�e �j�vr.
S�#$9T-F:c�)��{��W�]�jt����SBdŽ���������j�(�@R�W�Ō����x��P��S�r�`�y�zx̬���
ѻ����F-�|�Of0�A�� �,�H��_�7�%]܈{|�b�&���ʇQu99b�*�Tr骎V9|k�_.N#Vb��hL��Z�{Q�����)�&��P%^Y���c��eA	B�RN��e�FELe��3)�fDI� ������Ҫ�os�5��1�A�Yk*bf{�*��4.���\�е��I�DJ���#2�Z��ȻN��"�z��$��#�x�/�
��u9�2I��S[̫��汌�.PD���qs��d�&����Pt�L�ǜ�ȣ�L�=�������<(��&.\D���PI�LT�<���Q�[�W��'�Č��1n���+1LTeT@���ɀ�	�$a�w���\K�L�UI���H3J)F�/*o*��-�]T�W1n_�:����rl��X�Xr*�Iȋ�wb��f:�d�c�������UJn���.�>H����#,��T\<*�!U��0&�Ud���D��
Q��,]�	�J����L�S�2_.�o�^����#�Y(�D��2��1/�������B�ٴ2�\�Ž̧�D��FUS��nս����Ԙ�sbMM̄`��B���(�����9Riࠞ�T)Y1Q�tb�����n��aM�)M�	��Z˙w�D�F=ILd	�&�JyS��7	�V�Y�ǥR^`**-��(RF������%UW���e�.�Ip�3�9���eD�����Ne�ɁE�Rqr"�ɑV&��*�����p��y	���˘���o"b\�Aw�{�Tړ7Ouu�%�.�|���P���$�S�	����^�E��&f/؃8��z����4��!A`�w|�5���WT)�c�`��0���
�b��<�x�ÈM���R���>�d�Yz������>�S��;Hq�$��j�#� F �!.�2�fZ�a���j� .�R�Y�Uhh �%��]� ��St�  Ղ� �Z�j4VT��� � ��w�� @J�I1v* %���$J��SnE��Acwv�B@�E��!vD�@e�@��	  XЀEܠ]��@����)1K��Q .�(j�f�����M9!�fAAdlX�@���4H A	��]���L��i@@p@p�R"
B��Eʸ�v/qX�@��l������KG���?S�(P?'Hf���՗���>	����z����ȴ���:����s���㿟w��m9�yq6�zi��w��7��1��~~�}��c����絁�C�ҒO�,d!!Č(S�6	T�ۺ�$�������'�?�z��C���65&��+n��\�%�4��1i���K�ʗ��(�ƚ�;C7�!U�����H�@���;kB�\��t	�f#��j�h�Q��	s�5����-F9�����b[�4����5�}`��)f���6�����څ������8R�":�M����f���s[k�r��lK+��[ �T��Pu���MK.�	���6��L�MX*F�kc����))�UΕ�*����[��Ae�]�-��ͭ.�!Ц�[cD����]�eq����q�j�F���	��cfUQ��.�4�Ƙ1�.���6tJ�a�3H��b�\:��#ܘV�Y�������DMkJX#@�R6k�أ�3���Ҙ�<ٚh�ZE�F�l$��c�(]5���m%���'	�`���s��_�q�Au�3l"�pW
׋l��u�6�4��Li��Z,���ghm�]j[��f�/1���b�6�t҈0�jL�X��Z�X��JXg���88#��q.�n(0R�&J7p-͢0Ы��U+�m����퀊$�O;�oh^�m�V#r<�LЫ�� cGZ�v1�jHg��YZ2�#؈Yl���0Px�G�#��/�v�k�wp1��DevbV�(������	n��l�F��k��tɰr��e�Xm�V�x31���l���h��av� 8��7f�ޢWE�`��f�b��hA�ay����:��@%L����Am&h�	c�H��e.�c@��)��w%֚.�t�#[�`X�Z��%
���hM,1ί#ͩ)(%���k\�K)V�v��u���f#c-�t�Knd��S �; gf��kf�L�p�5�Pf��Aqc��e��3W�H�ik�5�`��7�v��b��1��X �mtr�L4n�n+f���	�K��3Άn����%��G�:�f��nf���V��D���j=IaJ,2�keb"F�b�\D�T5ĮB6�Њ汎��3M���Pwg��Ţ˝0J� �Z����kN�R���Q4"��F�6f����b�4y]a5&[.HL����1a�/_�ߓ������}�|����@ B3|����9{���!DC�g./�]�}���ݼ�@= �/����g/������=��j�qẄ́�{��?�޼��~�?`>�Ua阺k����F�m��S3�ט��{�8�:x���'l���Q�2(��C3Z�7�Aκ�S�p3�p��ϫ ��u���"���薞����t�P��<�l�D�'ŔoON7>Zt!�t��;��<���oZb�m!��m�u�T�M�y����|��1W��DB�Me'�e��W�O.���Y�R�����N�Ya(N,�����)�◠un;T�8�/6�IBw��͞m�?�7�՚Y/oI�)�3JI��JKY��x��nОk/mͽÒ����ټ��-�^�>B��5��<�,e"�bF� $�g���6���o^i/���&�XN�>k��w	�e�����1U�QA�!�x������6]��o|�Ow�w���>���t���[+����3D�=�nbI���2i��o.<e�$�r��,x���^�h�6B52,^4��%ċy�E��бB�C��� Bi(A.���S7c�O��ml�y��ʯL��ｙ�Ͼ��e�ď�>:�;q|�f{K*������cӷm��/&���;�LN��.�{�������,��ʐ�>��E[ς2�=�L�&$㬁X�<gt�`��d��A�hpJ� ;�Q��4�Xk1N����s�_4��wkg��l��b��̓�d����|a� q>��)m$$�����a'R���ow1;w�ݴ������K���7Yh^����>��xWo[WI"��<Y�F+x\�ӈy0M�T��1N�I� ��$%H�r���2,(������9{�T��"T®�O0Y�ڗwo}�i��Yo��f)F��ֳW��|�N�k��<Aq/΋/��v�O<�פ��j�2ٌua@����7o�D�E�|t�Vd��ЕӁ5h��Ż��w���v��+e���nxb{9=���:���0gyv�NB�AQ0���kr\V�rq9�s:�1����3���Qۖi��%�@of��K�g�bD�9T�f!������ X\�;�:`�!n �7�&�Y23&0Xq��;�Û�8�S7��p)1$�Yގ��1�8�}N��#���c���sHs��'n��2ȗR�q��3���C]B�����Y�%C;3�I��[1"t�IJٵ���lF4��W�Ús�/j��� LI 2Ww�ޮ�>'������������r�U	a�@2� MY"�HB-.�Z"�E!V)ݛ��A Z& Au��~Tے].�z���$��yiݏ��~��k4=X�UYP�YP5 5R�	����* ( �,��UV�6l�zmt�AdiWr$��(ݱL��Зa,��82?@94�P��!
KGDi��غŶ��F�a�5��wFw��.���ʶ�XmC����5�nv&�5��*��ٮ%�5��$�*`�N[���:5n�\Y� @��J�,,nȅ��:b���[m����RQ�PJCvB��&q�Z	H%K�pm6i�ʁU�4 �x͓6�шP���4��F�/cm1M-�*�gP.��V56���V�Ң��:��G�f]�H��'τ�����6�J�EiF�Z)���rJrMIt���РrA͒���Ia�o)�����������ߕX E�ٳ@L��+8��{[9X`���M9f�9��i��]��wlp�ܶ��h4��)�3f���#5�Сhu�k]��n�s���]d�Iˋ�	�[�rL;��"�0�4�ކ���s/qۛb�ϚX�N1&}���^p�נS���`ഷ�z������ԗ�{�v�p�H2�� 3:O��w��,���6�b��"a9�P9�&@�`����	�i�x7na� �j��L�[ki�-�>�
� �9������;�b��>������56��>�h V@b���_3�H��N,����W�CM����bk<@0V㍶a;>oP�� ��ي~w�j�T�3*7nݑ9>�oX��[Km���l�j�CPj�I�z6��GoS��#.ɽp��ƽ�ilk�6����3��0�%�J �B�I�ؼ<����;��`iaM�`�@;�q�f�`�ۘ�=^gi����S��o޾g޷ˀ$
"�	G���&'y�B�أbHX�٢���pB�@ER����]���-����.�e������=��B-ŷO5�R�ی:��k^�N�A�T�s�'xt�RQ��� ��m��nx>����1omk�S��ӺH���yܓ�}���U�|_�˙	n`bn���r��K��p�7�	,tn۽Oy��@�l��r/p]��� &��>Pm�� ;o)��8i�7�P���-��߿gk�KӲvgi�r�.v"�΢ z=l�	ݨ^��ig`!����-S��S�P%��=v2������ѭ��<��SxmҏX5��}ٙLș!\ʲ��ؖ5���׾:O]�pt�÷��z��?������bޝ��Y�:�в�[��V�ɘ^t i�O��q�5�=[5l`S̨Q���/b���%(�p5�=a�F�ǣ�մ�&��\7�� �4Ƶ�S�8k�����S�9_d��{[�g��I����ϝq$� ��ȓf�}uA�0�|Ͻy�#RKA�C�3�dϔ(��H9-��Jm
z�i��f�D�!(i.��Y��[U1�t�%�H�y��͘MH��
ő�X~��>q���L��v�[0	�T3�����b���'��-�v�f�����^K�l��g{�9�2��-.M�p�;�=s'M>�0��j���*\�+��P�͕s�7���]o[מ����:I� �
 a)a�UoO�L6�����@n���0��� O��
�-��
fy�P�;�k��$�L�9�M���}�|�zq��=.̛��p5���H%�~`ӓ����O�:M)gF�Ω�G�c����^)$��(��0*`G�n�T�o9"��K�"c�8���U/"�c����>	Ir�K�	54rf�,/bc>xzK��8�u�i��ϫ��fU��3C�Oa9{xŊ~��P�q5�����e��&�K��!��|>K�h��W8i���ԁ�qC�!�����"�4���Aߜ�i����<;���R"�QL�g��X�x�M����;�<p+ ��=}��E���,�ɼF�u�D���$��A��a���0�	<*��F�l��y�8�@k�	�%|$ql2�E���a�f,M�m`|G- ��x'�_�kc�p��7��I�<�����}!��ۏ��q�L��ú�(��\�'��
 p�cJ����L(�Ұ�:[���qP���f�fV��<�&��i 6gK4�~V��A}���}��XBƀcy�˔oTm�.�7UR.�7��"�P���g5�������3���A�	e�.1��j�lHj�Z��bY�H���ӠC��kr�v�ˠ� �D<<;W I[�g�}�C��9��f����ow�	��kmXp�A׳-�bG�-o�I�υ����N����Ǟ�;���2)+��C�f`�4��	���ʇ�n@Ȑ�rމt��d�f�H�d��_�N�6�6dz5�M� [���4���#�x^;qE\w4���s�w�/Èw�%<*oc�p�1~f�""t�cd9�4�\HE:��GP�H���/�Ѓ���oz�2�-Ly�d�;I8��|l�y)�>b ��c�]/�p1���f�X+ir���'�v�Hy|�v>�5�������<�8�4�����65
,���]�&۔�4��$jPvq^���;�kē� `���M۽��ư���5	���<�-�cZ�\WV.]޽�hw����~ϦY�6V���X�L��S���H�GoT)�e@ k��eg)s�6k��'����"!���DD�D���U<�l[zgϞ�|����]ԯ���]��c`g&.G̛#]��]k6�F �l�-���'���Ffn���<`��]K��LXЦY����O�}1 �cK�Kv0Tt���xi���:Z�xc�u���Hk�,�hlS����#�`��딼�|��~o�wx���3Mn"��p�xv�.F�0:m�<�:�N=ǈ���_P��,Ѐ"L60L훸�OH�dq��L|�l�`�Z���Wt8�r���,��o�'o$�vI��C6�H`I�'�$��@
.7o��p����Dý��4��&H�C��v���I���1�R�美A�l!�?sҟd����l��7\���4ណ�84���xP����Ge-�7�<����7�=��w4x{�dw�+-�Q��Z��ԷlX�@@x�}7z�m���e���dѾ���S���OQ-�xZű��s�iw^؂��V4D�����������| h��d<��PX7-�C�v���&�������y�%��ke�H����@�8з�{k: 0IL
�t�ZP���	�$@� ���1$bf�"�5@( 	� J�wϛ{0^����B�<�~���p���@��眊�3FW���ǚw��~�����}�1U�`�}e�$DS�����xȱ�9QX^dH�Q*0 y�z�0�Z��/�o1�=�j3��^xڐ�/a�W�v�3�=S3�ʍ����y=g��B�*��_��g�<g��Ȯ�^��|�|κ��7������� B@�E颀�Q) ��D(DL2��،75V,b�F;O����B'�^�U���.��W��sz�V�W ;��Rݒ��K�6��H����l��l��](�gB<�A�XQ.�B�E���in���fRi��l�&�V9RR�s�
JbQ5-0͘���M�h�at�9�(kaKJ����pث3X��"`���V�&�.6j������P���u�Z۶`Cl�ڛR�K���hWA����3��\�d1��j�ahefc�+�:����R}�>�2��r�u_�_9���Ơ��FŢ//�ٶ�*��ϲ�gu1�b��&�h�3]5����HI�JC�V�-����Y6e_��чq�y,V]J��
%�3��S�����ߖ����7�����́>-��Cbd��8� M�\h��]{�� �ǘ�ܘH�8q˷�-���'��� �<�w���Km�9[��wB��������ih�>�,�"������w�>�:�%�SWS��m2��me�I6���_+:`Rl5�y�l�2wu^U�W�U��y�-3Z1���D"Ix��"�H��a���r;4cla�su�:"t�A������� Y��і�Lkx�g���X#��hA��W��'�$[�m8z�4w�2w����Xf+�����s�4�ou���*��E���%w�Hn"M�Z��Z�8m̀�:o�:^~����F<P����|y��#���D;kKY��30";��"��\sV���t�H{�'���~�Ν<�4�2��� qXXX��׵�'�D0p�o{�Kqlke�Cc�U{�H��""�	�fH��b{Q����*���A�tZ� J�OI�n�Ʃ�q�xM�6	��h�:���
$�TkqҚipz��B�<���,705�[*�U�E\�H��]�wx��"�5����[N1��[�WO $����0��@� i䧞lPXi 6��*��� ԇ w����vw�����\2�FW	C��ۊػo_8�.;��]���EfL�G�9��W�'�X�֢aoC�-`s*���
\������"�`�2UP*%�')LAO(O�Ș��b@�2Ǉx;#d{�{,�# �;y�N��=$�afU��<A�e�a���1N)ä
<h�x�ރ#O��k��s��A"'Iʈ����wP�AJ!���ӬY��i���8Z���[o�Ķ�V�Ka�c�OK��h:��z.��=����؁���4& �~v�:Ї�g����ffcr.��a�y��6}�NVL7k��A$Ia�GtV��\��(��D���e0��l��^{2ÎU�sۮ�W��g�@(A�������V;�B�����"��y��/�AQ �Y$o�κ�^u{��7Q.&���Ml��;����v� </��ݙjhb��K��,�?]����^5���@��$ �D8�b�@7ʎ�)+��;�-dA��]fu�P�k"E��ܲ��j��=�����4��`��M��~O�Ϝ۽�,uY�l38LB�<Q q�݁#Em?	a� L?VUq�ǧ��3�:,c���y�}q5�Yfv;�Ƹ�'���Bαh}$6��I[-6@��c�Ȁ�$;��^wP�;�(���.�6��l]�����7�!� &�W><�"ZP�v;R��WU:"jD<�q	��z�ס�M�5aE_�<�竿x� �h{ ��ժ}1r^���[�4�/l	!�$�������_��N�v�Q6\97�n=jAqC^m�����Z�N<�/T��N)�eR/5�O���5h��>V��-g������Q����Br���
>��+�yA]�ӣ�jf=+=d��r��C,�q�:@��TUQE,�U!HPDRA�A@��H4�H�/HZDр$�NགྷΗs���_fx��ka{,<��?�N��E%+{�1S2"��F��Hl�=I�ǜ����$ǳ<q�tً
�>��D
cLo�;0G��`jj#Nsx�s� �R�XNt�Ķ��y�1L`lϿ��/鴝�cqC-h�+��DD=(�Æ��27�VŴ@�F�\	n4oT¸��ljcXb�Or�Q-�`���a�6_�DDD��aG㳉�n]�Ϝ���=���6:�u�z��� ��(B~��뱻5�%V�L$GR�ƍ�K`�,���t�封e�(���!+�1H�fH�^d�j���;6�#r���v>d�%��6�s��2�4�p�t�[�:XA��ـ,7��!�lpD�-�-y�{!�H[�,�XH��@S3B.�w�'0@Q�W�Ȅ�N�}��+��[��q'� ��zN�VS�c"!�iM����k�,@�<d�u[�
:Y��}y�e��IZ}���݄��'5��`�W]lr�Ϸ�sﹽ^�{Us�Y���bgF�?��4Z|0��bV'
7���}|HA�3�Z�S-c�� _A�o�x��Mm�1B^�w�2�j�c0� �U|��<:�`x	���=̚�0Zt�U�:\ܦY��� ��C��w��8�T���:����zNpmt��8���m��{�)s˄��j�n8E�H���B��d����!�S��K\�Z[����g��=����� ��wd�9��ÓY�~1 "�b�X��������71�g޺���:���y��vT�` �b�ћ��86aG0ͭ$V�l�ܰ��[a5���n���o)9hiY1��Pc6�SF+pe�<[s=��>����o=��8���L�<� U�6@�cxͰ<h1mc$8�&�p��GL��|��{|��"^CYyf�ȔO�����B�:��i�Kip=۪ h���y�ɧ��8[�n�[NF�sm̭�mpx��T� ��>���KgS'�ܗ^�ϋ��(df�vm�LC� 'xv�bH�۬��%� vHZ�&W?8y��LP�E�a\��9�����&3��z��Z�!Dx�E���x-<�`�ٟCw<BJ�Dwn�a�]��ݼ��I�0�=?1d�h�~m��51�I6�7\�ƍ�Ӈ���JXqX�x��۩�+2-�>-� 0ۅ��&/�<�϶ygO�G��{���` G2�f^D� ��7��ｐ'�^A8�2����q-�Q�
b���O�I=+KI�&Ho�x�+$ c�4���\Zၫ�%F�@%R���s�5a�+�s��	��s��dD	��P���s��'9� j4���9 =I/��g������}/?&јuW�>�R���P�/��"�{���&�Ԋ0
c�&(��y'�*g��OoA<^F����)���R�W	躳Q�T3�k[�+�Mkֱ�*t��g�w�Jl�s�o^9��Uwj����[�FDT�GԎz#�EMӪ�)��>_v���tw|�����j�2,�JH
BKE�l0��)�A
�5tP "�/�*�."�A�@1K22����e�}K���E"�6c-fQm6g%�� r���tH1�9�P�,]�!i����Q� �-�J���\���G�@X��i[�괥B�4���Xm�J�a4q%�yc�m�mPe��\�l�l��I�h3XZgZm�c�Pɚ�b�\�d�n�ͥ��],����p�V�X��0v˒����	��jk�y��ŰC k֚֫��2a��Z:��T��xh�^�w�i��X�
(
LfM)����hh
(b���)E5A4%�	�4.C�D8Hi�* �B�=���̎dW"�^y�� �j.Tm��E��kW�b��fwr����Sbf�\��f�$�ݤ
^P�i[4�nl��5�`�N��w(�ח�vWk�t�,@���<L3CU���e�~|���i	��m� �\zØ���Qf�}�g�� �����Y���� �I[�����1� 쓱q��Sh����@D��W��L��z{{X`�nn�x�Cg�E<��¡]3x0���"�3^���Ǎ�ɶ�����@� �k/�X�<�,�GM�!�>ʯv?(�fɳX�#���zŵ�6F���ی��a����\'�@�b*cjĨs|+k66��� ��f9:Z׀}q.F����Ą�����U�e�c �W+���r4��3�R�y��(i���-�K>�~bH�7:�/�l��'Oa#r^�q�\t�n���C3{[-��sʿ��>����^��d��2�nj^������y�$������߯ˤ�X�,|d��|�rÍ �k!7��O�k;[R�I�.[�H4���, �3]���������t�P I�#���ŝ9��<7�Г⌀" �B&"ah����ޭ��a-[u���jҢ�Ҵ	��8�Rcpݬ&�A�@�
����
	�6� L��5���h�������s��##���'���^n�ā>��w�d#-��	n2�Cg���;�/�(�yC88������[��|�*f]��C�/�@���<!D�,�d	��W<�)٣�j I����Xqa�x.��>�p'Ū��8@����~M%��6���兤W�_��y}]Nz��f�*e��Y�3���O
����&'{=���砷_���1�1m,�p�X�g�M�AA�`{N�G[��7�:�������!rm��\x��:.�Eq����y��f@���݂032!�C�<>�8n�PC�]�/�60��@��e�al`	>4@�����������3����s�m�ӡ�� W��i�${E���R����i��O�rO����>��6U�9D�0�-#ꖪ��oG�2af~��m!��4�ś`x����`�F�\��KQa��;mo;4�l���<�|� @�����V�٣3��s�J�rg��;���Ϳ~�\���U���n�P���-���#,ɵõ5x�x ie��A�[,�ڨ�c�.G)����PŨ`\���w�y�l��~�rs�ac��:x��C�����[�X#K	)�zݚm���#��>�K�.Y��-d.n��fD"�L��rTDDR"b`Ϙ��1h��ݗx���=]C`e���0��=� 	�1��yoB� q��`�����"|���|��.�����r]��Q��Rt�ӈO+�m2_��w��x>b���<m�鴰s�9�<���L�4�f�=�r���=�خ�%�b<�_�'=��`��a�j�.ǉ��th�WT��M�v>03�ʀb�Ҝ�'�D�x�&v}���k]�N�[�P�<����>x�шڰnu��Z��+#H�"n�y5����@yq���utK�[q~�^;3�X��)Ɣ�rQ�u�:D��If$d*�����(ihj��
�ZR�J��*H�V��i
V*@�"���
� ���*
ZY��ji��)\1�N�5$��R`,���=zu��\�C��p'Ź�6[�s�b� �S
�'-�)�t�-1��awC��-�I��!y�y����<������Qm-O�G{�0�!Ǝ�]BEW�� ο����-g��8"�U5PhE(��	D$��r�.H���mb)�����}X��N�o_t�ca&¼.�S�4�jM�}��w��ꮼ���>J瞢$
I��Eb�m� �!�'�������~w�]��w��E �,�s����.^s£.��͛KYhn�Y���L� ��1�%�f�, ��V%L"� \�J"��:|[<���*�O`Y�����눉�U��l>�Q"ǂ��]� @枞@O���z��.�"2@-�+2\Q�P�O�G���x�W��O�\o���(�R�4FLW*�ii:wä���0{@����k�Ao4wI���K8/>�yw�ߧ�>�{��7j��a��ȹ û�a\�
 ����^�{�-F��3�Z���� ��:s�x���U>��~|�Z�o	��D7�#ܫ��ee��� �@H�-��DBf��K�7���������y���P|���	����x��gͦ��@"�����v��1��L� �V���yl��d;��"�N�.��!:x!�xb
)�i� �1��x�C�:[�4ބ�"�@�X��wy�@�Ck<`	�b`����4~��wۀ��,5b2��^Xש�l��@�3r����"""!�PA@Z�x���3[����P�X]5�,i��U+aKB�m.��%�H\ؘul,�PV2Z.qh�6��\CÁ��#	�L�+D�=���QZ��p���, 1���Ys��]�kɨ��D	�~��0��gF���貪�[�0r��`�TN�v��`Lw� ��U{[��$�A��T�����y�ip"��$�yKW+tux��.up�nL:�e�muĵ�����ߚOt;>�߆=�z4&�����v����z�^5�&��齇ͧ�� FL	���o�5����%�㝹C�:afߍX#��:N�@k�yک����ſqb(���e�~Nt�T<-g&�������w����9Y��	gQ�Us(&JcH.F7�P9y�6���'F7�ప�d�5�e⬯i2��0�)�ҩ-L9PD�bK���:�"����x��2(y�/[�Z��?~��K�ޢe�c0������q��g�@AvZ�!�,|Ψ�|�o<��e� ���e�rT��\��Vg��;N���\�/��g��ҍXa[���K�DX� j�!cZ���@��i�Dլh�� DE�&RɉpK�6� m�|�����޽�m�߈�ί�˳�՟c]�[��At�H*�V��Uط�/[Ӣ�*����N� ᒂ��dQs$&8Nz'�^��c�]������<��>���Rr�����dL|t�n��H�����^��R����A�x�U^��P�"�ˣ�R��X�S ǋ�>����W.�*�S̽i>Vb�T���X�lk��ﺓ.F,lZZ� ��j����VHiH	L&]��2D����h����p
1V5�EP?w���æ�+ǔ�f�l��cYWP���۵#��2��MH�������u�<�@ŬIiG<�k��]��u3��q���ׄ-3�\kmeD0�k.��l�	��^\�,�&΂l�3M)V�mt�l6nyis)��;�:�\õs6b��ƙ���ftc�R�H�QL�%[��[
� �[��oa�����ie
�"���D�����gcT5�B9����)�IJN�R@�OD�wN�Jw����=}7�U�W`��M̹����1)�DId�w7����ɒ���َ�0A��V\�k��mt��bKN�6�̳R����r��D�b;Ɍ�):�O�:Ї�b3��I�O�Sm� �x#��
���Lu���v�-������2���R��LW��#�������r*�mu¦%���2�� A��=��� �M�����%O;�
�@�#���s�-��� Y�ku��c���i�H
&�t ��2��G7vP���z�����!���xb�B�-G��-�l�	�>�kga�n}ݿ)f��iq��7K�*��w8�a:��M1nc����<���R�͵â� %��8�]��$��	<	��k-zc�w\DKx�>-g�<�}qM�lel@�:睥_���,���f�$D�q�{���3�W�j��h��!�[˶����Tn6�,ʉUwO>NI=���7�Xv2t���[�<��a~B��0U�� 4�q���[��O1a�Ϸ��g��A�@�q���,���r.���>C�4DDE��!*��ZL�����.�A�����#���"�T!x(гG<]�if�oAp�;lrI��r,��*�2P�� ��(���a����ݶ��j`�dނ&���e�ّں�����xv��#N�ݜ�vw�)D<r�a��hە;'����%���A2��t�p�ڲ�\!�W˯)G���30`�#��h㞸��(�<�X[f��R�t�0���J��K��X���?�{�w��e�Bl*�]U9ZZ�
�xF���Y��4�]����1�M��(�ûtU�niN� `��%ʺq<ܺ�x�:� !�6�~��=����uU��m��E�d�5�;��m�3kK!����<��t�b�Z���ʀ!����O�a�(L�����*T�3��0~��!��q������g���Lk�� �˳K�C�6�hTY�-~R��t����z���kc��u�E(�a��9�+�׵�|ڙ�M���f���L��n^��%�>���7��u>w~w���B���zۼ�V�ۘJp���ֺ6aq606�P%�@X@�JC�b��Il'�;����y
96b"ds���sϔ������z�w���m3����h�N��0�cͱn2t� kI0����cbSx�>�ʆ5��<��⊔�i�������aD;޷a<�8�HO��yk�[��J��^����u�'��u싐�4lrk"[��O2/��c�(B�kw[�yӁ��E���?Ib�Ӭ��&�.��`�DQ�`K�A�a,|���@�F��R;�d,]��/o-�V 3i�P�է�=�~�'�Ǌ���"Ϳ�}3~�jj/<mT7cי&;ݚ�z�S躥�g���,���d�	�����b|�L�qRP�z��y��T�D�K��{��L�zk-��'��ʃ*�h@���K} ��Z��VSᗔ��7�eI]�1�`弋��p�Q��]5=k��T7֦�����_N����Q礩(|37TZ�*���:�6�yo��	�]�G�Oq-�Q�1��hB+�5S5D*�����Y`ms~;�&=��<�}p���y c-�|�:ZH�E����x	��`Yn�5��>�I\:�Y�pjmPM�z s����S�U�0�0J��.��[�vv�g�\	mbxS��,�6��ў Q�,�$矪CpX�!�������8Buu��מ��hB��fo��˻�o��ξ^w�}�����; AU\�"�GjsL`u�2L�ٹ��F�G=��P�K-��K��M��[2��q�y������]�s������!�+/�F�~��]9��3T�����ʋh�� X�,��d��Mw�p&m`l��B,� T����	Ρ�(!ϱ�Y��ˉz�s�p���]J��S�#Y�3��v:Xy��O3a0F �կ�:ZH�LXo1�v��Y�u���~y�ޒ�k4�hY�"s,8���m;:����k;��Y�%�ZzPF��x�u���"�7D�X�@�6 ���b�^�i����y埿?����B�w4*�J.LS���!��<BńH'��3����7!P,2��H=<�gM����C�܀Lt��ب� ch�c3J���,�c��< � `3"d@1���쀴��7ϗ������}����8l��殞B[K9�j��<T����!��<o��N��(i�j<�" ����y2�ɞ�fϬ������y�%O�X`O�y��ZSf�����gi���%�-�[-�) [i�KB��z��&(fUM��曯[%g�����.�@r�ੁv��p$l
N���,D��x�ko!G�L-~p%�*-��߀���6
Zlˎ�Р@I(�!��$C�x.<BRi���f�4��PG��%vB�.�D���1��>i Ao4Ϻ� e�4GF��XI��p��JG`[@6[��̰��I;�Ø	<;�r0��M3���WWD���6��-m���4��GX�����ċ�ʹ�q�-�Ě*z[ő���p#��=��
f����������#Wa�c8�i��'l���,�>���ƈl��e.Ǧ`�!��%�t8�̤�����k�w:n�[ũn�!�^�Ha㠶�$�4u����2�.���g�¹'O��:z�� �I��0�o���4V�)� KnMe�i�����F?q���;���W˯vy����]�Vܩ{�%���r�
 @D@X� �E�,j��,h@��C��)���5d
Z1,��J��C�:E�#Q	�1�Baӌ!X�m�EB񘈉���C�zS8����c��C�D��3tC�a���S��9�h��ޕ/S�w���ڀ�<=3b̌8.5��d>TO��Ǯ^Ӫ��!�����<�5�x@�T�YT��y�3��M�Sr�9wR���Yy�W�=�F�	����ǉǙC*#3諌��I%�s耀�5`EH���m�E@B� "ha�jX���#�K�j Wv؟
�0`�,�� F�Q��6�RۛW�Q�v�p���Ll���X�;M2g�.�hGC�qj�с4��]�c��]��1.��hVк[�Q�YhMv�kVX�-X\R\�D6ɴŅ�u6�[v����o-('CrY���mXL01*K,��0%&����#h9$έ	\E٥"�	�*sdA�Yk� G�1����l��s�J�6+b<�]�F�j��f5t�7�|��H�� Q�(�h9ؗ<���*��q�}�}O���U��+("�3<���r_T�^<V;dFA-3��qUkd�떥���[�X�7[(��ZP�sv݉��dW�c*V�b2��J,��xf����!�����=)L�>b�/0�U�t���0��w;�K^�g���A�O�Kik�/�r4L�mvR�M�V��o�f$���zc��|�:@z�BHBG6brn'٬4q��c�V��PL8׈Hq0���l�1����}���7����@����M��Յv�iz:O^>x�v���&
�q8zJj:Dc$�^��8 ��,t��P��d�y�}dF
=��|�- �o3��S�q��cG~��<��^w���e��������9��|�Kp��r7��-�8�&:+WJ��&<��0�OO)��5��	�|�cb&|hK��Wݶ�ں������"@�<��Ű�Ȟ���û��	˨��(J<D[idu���|b�/��;��1��ߞt����b��L+�p�mɤ��-y�{!�8д�����0�P�Wr���������ߏ����o�|��*����(F+�Y��J���R�)��Kr��02�nD��Ҝf�K, c���P\��VM�X��z�ݮ�2���*��1��D��L��6�E�9]��2����`p� k�r8��
���G{s��H��h{;��с��ȃ�"b-e�K\���7>����ޟ��=� ���||(��O���j"�v�z��]k����'za�t޶�<�4Z��~y�_�|�����7�Af��X��"`�"�����`��[���7%�F�*�j�R��x4��a8�c�;f�'�m�;Kd*���z��'�d��{�c����C�+ja&1�/�}���+��]�^�f�z��U�Uû��n��lo⏮��`�\x٧��^��������<#$���񎴂�	�5ז����}s�F�z%���4h�!-���OOA���c�@jw�4��N�I��i�v�h�@)@����ff��u����WÞ^��>u����7�Щ-����y�6�J��)�vs4]61���	I)k��Ĵ�[m���%c�,�eU
ܕj"�JrL����'��1�WT^��6@bCH�UץX���i<m��XE��8��u_>�5m�f�y����lw��X�#����P@���]�e.�7���������9��7�� ¾��=�m�y���ZBv�m��a�`����r��5�2�&Fʙ.�K�t"LCH�&&GWx Nz�yv>���Y��ܫ���}�}Q��"Q�]�g�fx�O���6�-W�;����������=�vUҦ��bը���{/d1"ɴ}�1W��}���y�Bly枒)a��
=R���"}���1�V�$�=�Y�QH��1N*��7')ay�@�������򸧹�����EV�g�T{")��i�F�,�V�OeN<�t�$����+�PBe��9�ؑ�\�(����
�b+c3�9Cj��4��*' ��(h)+3"&��� ���a��bf$�i�	&	��X�j�	�Be�K#$d�I�)a��I �d�q��X�d��B	�q!�`�&H�	 �"&X� �3&d�h'3h�����
J� �(2���]�5ӏnQ.�M�hZ���σ�M�����L�<E�`�iḓ�7���}���ܩ������ۈ=���m�l���Oʬ0�#+�t�> �.����E�͉G�s�}t�@�wB�����z���`����qp�R�(͹�$��}�OP�����`^���	�������[�n)���C0����<0��^���X P�������L���y��ݾ�|���/\�[�s��ư�dF+�J�-+jL`�S����Z���Ye ;F�`iH@8��l�z���� �W�����D�M,�������ݐ�O-���[ld5h�Y�rl ����{f���pA䯅�'���?7�9˻޹i���T��n[��5��ѧ�w0g9�$���D5a؝d���h��%\2<&Z���O_,����x0=�q,��C����8վWt�W��Փ�˒�7�ļ�l������yXkf��R�}����4�<L+�v섔p���vk^E����"���eW�}o-��s07W[��a�&{��[3"e�1��s ��) ���rw�����\�[���P����6����50�:� ø��1q������wc�E: ʧ�x�Ӓ=�l*faDND@�qst°/�W��Iϳ����<�˩ �J�j�5p&��S�k�᧮���}���yײ�kD�bYZ�� $7'˙0�TP��>U�y/���&�B�!H�5-�2�Fܹѹ�W���q	XҒ�L�Kݴ.�&����7,qıՈFV<��;��.0u�������-��{����rzy��Jy�ٟ�P��ÿH�?z�E��еW�@��S&��;s[ih}�"�=�y��r�u֗)?=I;�!oC��`N�)�*�S��I���8}R�ٰ�@|���{h�۞�kG66�oO��>��� 
���J��l#t�;�#��OL+G�W.�½N[��<$E���x7YP,�^�z/���o&�A�~|f��^���[ma`v�I���2y� ;���e�&l������,�w���=~�az���I�O��TՃvߞ�l^���� ���"�+\�'{7~�:��ӑn�3O��q���fZC��]��w/�ID?-�5�l��k���y����#Q�o����p³Hb7ӝ����zw���}��	�O��0��i��H�&.5�UTUUUUR�z2`  ���Ο��ϡ:��H�gSM.�}Rp�MY�����N� ,28n#&I�!�kݘc�!�ti�o����p2��6�Q76�s\GXQ��13\hD��9蠘ȡ�K�� ��L 2t瀸`p�DP�)�D4% �-�PЀ�$��0�]S	 4��D�P4�Б��-�5����E�"a ;���@!��*���4�J���A������4����	i������� 9 !��"�H	���3 �$"����54��@���u�T0�pØz�<�C���F8!}2ǖ~$�3}�A�`3��G�<�S(0!��UU�+�D>@DT6}"&D����*)J�)@04!Q+�r� ���Z��h߀����s��9o��힀qq�`����������csn���	+��ƚ�č���jO��45/Ct0?���]-NF�v�6l��Ћ��@`h|��i�cP�����L����L��e_��X"*��M>���]���<������^�X}�{�i=$��?�Ǒ�*�������<N����?����v�j����( #��(	$DQO�p"d�M>�O�r��O�7��W���� :��a���
��:"}@� 4X�t�G�� '���#H�c�BuL�v��<�����~o�o��oץUW��?_����1��|>�d���>)��/9M�oz}�J�.]Ɗ�(}�B�b����饤���U4��W�!��'��@�0���NI�:MG������yr�ǟSd�O�3��LW�{j���h���}��^�}�ڱ驾�pR5.�3�gt!�_�>�ǮC�^u�읟iI�O��13@�0v릡�Sr��L��� 	VQ��GH(!bL�lPB�CB����
�*	@ЍHP�I�� C�	�KJ2�4� 4! ��" �C R� ��+BP��),��,��,����
�@�$���ı,�!C̒qSI�����	� A�	T1E`P�C$ L�G	Q8ˀa�M)�8�m���1��3+��������y��� O7�^w@⚭�O�ĉ��y�!�rS�(<�@H�K���8�����!�ww��h�<M���`{����׆���q"R��=��.����ؤ'��i����N.������s�}ϊ�>�J��{>_q�cC�������uS��{?0��ٰ� ���O��&]���7��M@���%E4�4�4��4��E%%%%%$�%%%-%%-$IM%%%%%%��444%��P����4��RP4�IBP�IIE����@P�RQIICICRP�RR���4�4��4���KKC2P�RP�RQ��4�4���II1II4����4��RP$�HRP�RDD��D4�4��4�4RR�-$4��4�IE%%BRL�3$IE$C�D���4��RRP̔0CICII1IICICP��1%RH�P�D4�%%%%$��P�R���RR��R�RP�R�HRP�P��R�RPP���44�4%��4�4�44����4�	ICIIE%%KKĔ4���RD%%$CIKE%)4�RP���$ICICICCIQC$�%%%P@@4�4��4�4��Ĕ���4��4��%%-%I�0CCD�ICIKICKCCD2RP����P�P�RRP����4��RP����D41%)IICPĔ�4��E1%I@D��4��$ICICICKIQII0�R�RP�D4D��4�3-	CRQRP�4��ICE-)CP�RP�RPRRD4�%%-%%)K%)@Ĵ44�RL�4�CĔ��R��P�P�$K1A2RP�D1-%��444�0KICE$�̔%%%%%CC@RRDP�P�P�RP���IICI�RR�D�R�D4�4�43%%%KKRP��$CICII��QIICCC�PĔ4QI@D41%%,IE%-�ICKICE,�CIKKICRDRD�4�ICIIE$�ICIICI�IP�D4��4�4RD�4�441IE%#D��1%��CC��4�0�@��̔443%4�%--%$IIICCIC@L�444��1%IAM1MUTTQS��15DM14PRDU�PPPD��(P��R@Hy���OOxa�8��4$�7A��ptdt=8 q8�@��9���1O�'��y!g�?<��~������Cۇg�w��j��^���O���|3ް���8�2}OC�7��<����#�#����~bh����}��W�=�f�׏�^�x������O1�=_W�U�=jm)�X�@���)j��}�y�Ƨ#���^>A�a�P��У�|����'ɀ��=�/�j�����M�q�#�*7�~�����m���s44�5��w�"��mG�1��C�`�{�?�jj.�p�&( #�f�^C�^�a$�قi�d;�e���D�;��l�+�OCQC�ˮ�x8"����|��	��#t#��ɸ�z|�n�o|�%H������蹠i�FY.��F�8��B'�����;�@�NC)��0��e�b��\�)��	����:���r�C�s��� ��yԫ�c:�dpEU@�&]�p·������'?��1��O���>TT��`�@?i ϸ�O�6��@��T~��jm��d�x{�q��Q�x���^��x{@�����q�������L��Oh< OZ}�����|���o�G��� 	~D�>(��%��������*�}�hrE�����������8/�O1�T����!�A��P� :�ı z�0G`>`8#�""�b��?M�;��rE�����a����g����6c���@��ۺ�(���`�����X �#9����<}P���x�"�fQp��p�XX�d���槿G��`�@�!��{����k�y��� H����/��0�|h9ǐp�B>�B���,5�U\?/�tiI���>ǉ��
��gk��᩵�{|H{�}�8�2Nu���`'!G��=� �)㹐�Fq��4�mՄ�Ą�8�^3|5�gN:��軁��W��BS� ��lL�t�Ë����NI��M���� 6@0�y�=�{{^���v{࢐�Z�v��L~��J���?� �a���O�j:��� �A$Џ÷��S��ù� �����'���16���L��S�_�x(iԍ�@r��
��|�!�'����sȧׇ�͠ip?��Y�}�p��̈́��>�=��A��X#$"� 7��(�����)� *