BZh91AY&SY���e߀ryg����������`�>�  ( :    �@      p  F�"�
��**�.�vB#���[p�������=���h�n�QӢ�n\�@N���X�)պ��CF�Ò��/y�У�3�(��9�q�@o@|����D�\衣���B�|y�_(��n_y���N�׹��o����\�h���W4(h8r�^�uy���ӫus@�ܹC�]�޸����W;�(��a�P��z(�3t⁣N�,��7� ���f�r��)V�(��@�X �              i�)R���&L���&����RF*Q�ɣ � hi���RDʤ�H2b ɦ��  i�T�S) `  �0 #F I�DM4@hh     4�&�z��z L��M14���L�L�yO2z�������'��s�� D��@���d���!$$'�@�]�Ӷݻ�+���ӵ��^N�V���v�o��?��>����~�<�?��h9�z?�/�>���<��v5�������:zu����������*��0 ��u4I۹!$��t�UO�cbf*��~^~�dHO��$�Ւ_�ǲ��３�3�0ԇA�������HC�o�S�0��$�^������A���I O���U$������ߛ�����z��g��a����������������=���?��9��w��t�
�aP�
	m�����5
��B�w�P�48���AH��nChT���0PX("�ACAA`�V۰���V
۠�݅am�r�B�PP�P��aXT
��aPPV�[�XT����+PPX(,

��{��AA`۠�*�B������V�AA`��\AA`���m��[��TAA`��P�V

�۰�	m�T+
�CN �XT
AaP�4��T-��v�B��
m�[m��(V
��WRWQ��(�E�q@,`T+
����¡�
°�3�t��m�XT+
�B��T0̨T-��{݅B��[t�B�Pơn��B��T+
��AV�hT+
�anA�
����T�m��AanB���Ь1�*��`��V
���A`���-��AaP�*���T*J�B��T�
	r����A.��շ{�Km��*�B��m�B��N�PXT+B��(+p-�Ь*�Ad��w%�sd��8� I�sd��B��
¡Pn(7>�a�0��)p*�1
0�[u
��Vj�aP�!PnIS4�*anaF�B�ơP�x�����!P���XV�V�T3-�����6��m
¡P�*�ӌ+
���*

�Bۭ ��PX("�B���
�aP�+
��P�,4��n�V
��TaP��P�1�t�w��B�PPXT*��1��`�PFІۘ�n�B�*�i-��t-�V�T1�*�B���V
ⅷAX(,*B�
�.ۘ��0�V�.`�XcP�V�*�`�p1�(V�*�V
۽i0��XVwx�'�NP��!�0��B�X%���P�*aP�Q�B�T��B��[�X"
�T+r"�B�*
�
¡XT*�p*P�VB��
�aP�6�Ha����B�XQ�B�B����,-�T�.��X(T��*��CmC�*��V
��p4�0�V
�aP�j
�hV��B�-B�XT+
!D+
!P��08C�8�{݅B�P���Q�T�(�am�{�P�-�[m���[�F
��Q�B�ۦ���
�)p*��CZ��!��P�)r�����m
��AdRcer�r�]ʻ���\�r_8�   �T��|ʜ�'9�/��?3�}�����=�Ifq��~�g>Μ������5���������0���'z�x�,�}:���oÇi�����C&	0Br�`�ؼ*t�ɃS��_U�Rr��N8��y���uBф ؋P��u���CN?�^����葊-4LI�p�<+�t��ʈ"�a3�2gL;���0^�ɜ1�d
�]d)�rnr�ͩƧ�?izo]Bz�}ӱ���=�<��}E��%L�H��5�>����T��O�q.�l�šT'6;�đm��Me�0(�7�N	Eã.P��`\Ș�{	*�{yȋ���o>T��R��:��N?�2D��I��*ꕛ�j�S��/'&�Q��]5H��+PC2V=)UK(U,{�&�M(Л�M�,��d��^G�Y��iR���qRO��:J<=SS3G����/"�<AȨ���SyN-=P�/*fNDd<���ˌ����.3(b�3s��u�=�����b1���R0H�����[�
d^d�\;њ	ڄ��!5��Ґ�8�A���3��K�M��+�D�|��.g&
q�U7N�"^��4\�K�b�j�Қ����LeB����le�	�l������D��{�zY ����2��e�lۓ�]���<��Ȋ��Ɋ�A�Ո��\� FHr�Z�t�S�N�j/.�����E<>)f��ɋz1/#idui���!TQ���=�-A�c���wR�z��
�*F����YQu4�w9Qs�*�[��"��ãyrAHY��!�oJ����**"�VM��˕��rr2�U�.���U�r�,�+@�\�F��D!HЙ�	r&���1!�TS�MU"�J��1	�P
�i�ʂ�D���>+
��:����9FfS�ẍ�RA#-�O�Ub��*k)c(�T��T���6(U��h]M�U����k��h,��)|<Fd=��)S��v��E�7�I1jF2�_*U��s,d��(���Wsi�c�\��B)C���R�@M;eMH��T��8/�F���{�y������xQS�L\�������D���yW���2ȷV2�,?�O��K*<b����Vb��ʨ��.�����H�"�*U�������
���9��f�,R�x^T�U��[���/j�bܾ�u)yT"*��/�=��Uܓ�j�ŗ��u(�|ǃ�	95/���ݫ�8]�|�tFY{���xUVB���`MT��ǧ��X*�/xX��"�
9S%E�ʧ�d�]����	Ř!�F;�&�Q�wte	&b_'/ݻ�ʄ/�heعy�{�O
�Ɍ���94(ݫ{ɛ�{��1v������W*�J	��Q�i�1��Rr���A=<�R�b��Ň�	Ǫ�y��R�7(W>��2�̉��z.���PMd�2�#"n1f�=`���J�(��TT[�*P��Ok9J�2���˔]R���3.g"s2%3�
ʉ�3
&eܜ��u��ʤ��D=��"�MfT*UM�/Sy.�!N�S���1!T
d�DĹ���2�h��&n���4K�]�t�M!NI̧�myuH�d���L�^	�q!��oO-8.i�� B�
�V��
k���S�R���7RaK��D��'�x34��˶1*�U��}��o����oc���!�� �o{7����*��� K��L�$ٖ���a(%ڂ$  K���` UZ $�`!Wr (n��� 5`��䖅(Z���1 B��*� �]���  ���L]��	cb��	�rTۑA,iX�ݭ� hl]�Q.�d�,m@ �4 w(k�)$cAm�LR��@�
�(�n�  &_��NAA7Y�PY&�,l2�Bn�d"��S3@e�B�� T������r� ]��V���[�V�_�>��ώ�|������g���������zuA2y�n�=<�ǳ�ٳ��׆�˶�y�n���://����#�	����z���!��0H�@y����:�$���_���O���׿�W���5�q[v�00ݠF�K���Xf�v!�Өu.�5�˖W��f����L[v ۍ�D F�o��R.SL:	��e��Ɍ�A��ب����֚�H��(k4�K�Hp׬�[����1�����,Y�c�[b�R�3Cjnc#�kG$�Jp��A6�R�1�短��]ې�T+bY]4�� �������y�)�ն&�U�Ը�
��T��L��35L$H�k�rA�ԛ�!1ɳ3Sq2Ch�[q6Z#r�o29��fL�v�[[H]����{�%Ҷj��[sZ�����]iM�0cV\�c�(l蕆�Xf�%&��H�u�BF�0���B9]][�ٖ��֔(�F���t�6�Ml.�>z`�)P�2�ԈE�X��:j�\9�`��K�-J�W��3��cۥ��j
sk-���{�ʦEa6���m�±0Vk��jB�Nɦ)eu A��=Nak�Ue����:5���{:���]4� �-ړ84r����b��]t����Vb�gwsn%֭�
P��F��a��FstJ�tM����D���wm���ʹj�nG��r�@)l�t6�,�(U�����94[&�LXњ����ۦR�Zv��T�z��tt`:�0�X���fercf
�-����v�+A�Yq[ysm2ܬ6�+X<��J��T76�a[��V�H�c/\�y0�66�R��Rix�H�,�������|�W�B]F7))�fd#5*L�Dm�������[�j�mZkF���8.V�GCiIB���jKLE3���jJD�	e#���2R�U�]�����Sft�ə���m�a���LDp쁝�]�c���Ե%n�n���Fj�]iƕ��	 �4K)QV�t���)a��l�6*ceT������hݢ⹕�[��Ti����6^2b:�n�@�SD��#m�6X��˶H�LCM��*nH�Z,2�keb"F�b�\D�T5ĮB6�Њ汉��.Kv`�׮�[���s0J� �Z���kN�R���5i,Yq5tGAͭ%�L�ERi��,K�:�B�gZ�_����n�{}���^���<$�Ē@��8��f�S����?������ Blz��;����'�Y ����۩�<|}�����/�<�ΐ���~�'��o�N���>�>���z||����&����w�j(q��Hfd=3$�8M�M� ��E�F���x��!F\ȣ\M9͵�7�A�4C`��2�f��É�>w�v�nkQC�oF���!���sa�I���OZ���t!�tB�ף�_��y��N�����t�EP9XI�8�z|����7��J��@��'��+��'���Y�g��3�g��:��	��z²	x���i�ĴC�#�e$K<�w��l�o�1�����{zO1Na��B��$a�(�/XO+^_r�[?/������,���xc�{.�'z�t�<1^�h�}3, �l�GM�-� &�_^Y���!Ħ�E;�p��J6U��b,�6��Ra�w�_[v��T6�o|�Ow�w���>���t���[)��[Re�j��71$ҋIC�4�} ��2�E�A�<^H{�B�LZ�ȱx�{x�-�e��B�
u
��a	������e*��kfB�;�l�y���W�f�����R��{�w��2��GΟ��N�_9ٞ�ʯ��4�1����{�ɻ������K��2�8F��ȗ� ∇�
�o>R�{<�PLI�Y��x2���/��Ɂx�����@w��%�i���2��q��s��N��Mf�:�^uw�d��&��N�8M�Ô"�On�RBE�����bqM-�s�\�L�IU*Is臟;��˜��
`�e�!����e	�s	ZF�*��Ř$b����=8�G����eJ-��Ě"	Q�A�T��)J
s"�JH{HѬ)C��PEK��%L*�K�w!EJ>/�>՞��@��#J\Y�CF��+���<���k�Hx��_΋/��|=���	��B&�������2�f��ݾ!�����Y���3�L[}��4vG��I|OF!�W�X��Ovs��<��v=�89�*@	��P�A��%�@�g!� .g�0q�8�i�`ua�'sH�
F2(��΀�6���C#"U��a4�:�ΘՁ�䘁�a� �ap�$��fzt����:S�#���o@i�o��\h�@�0���!K���g3=&�q�f�z �Ν-}r�ᓍd��L��g^2v��!�D�Y�%C92
�0��N��X�٘�3�I4�d��[5��ʬ��	>2HI D"���~�ēfC�{�h� O���������EA�l��&� VH���K�V��HD�
B7f�)D V��@Er�w"5U䭡��P,��2�/����&��}d	�H
��,j j��W(�T@P
YM&�� lٲ�� .���Ү�IQ�Ԯ��w��o'g%�����������j���w ��v�֍q4��p�R<��09���P�.��D&Ö��E����6���,
�)�\8�S�[Y��͠4e�0���-�B�`�ی��t���SLBƚ5"f�0��AAΒ��SUB$��v�pU�Y��1h���&m���Wh+hi]qIu��Y�^��ڔ��6$�m3�e�2,vXX�jKpL�����foyI�d���@��9`p�A[]m��Vص�T[s��p��4;�8ꠁ؆���S�0��ز���}��v/wO�|�;i�QA
ݛ4�˖�ܗ��X`���M���fl��4��c�ˠpF�-�l.Q��lLۤ/�f-+	�dPAC����LS��tR�P9�q�	���ӄ����~XoC��uO����ͱVg�,�'�>�Lޯ8lk�)��m�pZ[�a�odŀe�T�O	� ��Kn�IU���g|���I�$������b��"a9�P9�Y�@�`����	�i�x7na� �j��L�[ki�-���w:�>E���rs�x�5�����5C����M�!��O�����?��ƽ��A��K��̐K���{�4�[���L�&��n8�f�����I뜸�zƫ�uJ#2�v�)J��7�
��-����v6z�y��5b$�V�^أ�
7�Ȍ��d޸TZc^��4�5�`m������BMv�i���r�ߏ�\���r��^�4���0`�׸�M3z�x��P�3�4��mָaV��X�O�DDD@(E �w��͗n}ɼ��'N���.g�뿾O�y^NPH�@X!�cj5M�nWqt#.�s��7���A�@Z+g�X���-��iZ��8-�X�Q��f�۪�Ev�W��OR}}���v��ʶ�7���>�oS�ֻ50���;��+m������k��8$�"�Q����h�*��Y������Í��G|��=��`��1 �^�.� ٛg�C
�~r@m�=��0�j�٥�ӓ�$ŀe�	
	�Qь�^����*��n��w��r����J����N�	O�@�ǈ������&�;F�FLF���aM�=�J=`ׯ!�|o�s���쎭��dG�^CbW��
f󃦶�l#���O��oS�����chQ{��xYx+^�d�/�D"|TӍ��h�٨`��eB� 5�Z�canʒ|��z�����{z;m[Noz���zZ�
�A,k^U0��������;��NWru��=���V Q
!�D@�Kgθ�\�N��I�S�����r�O��^@�HԒ�B",W[0�uT�Q��vı�j[	��>P�	�b#fף&	�.إ�Ӥ�d��9͘MH��
ő�X�=���	��;xY���*�c���ѱL�~�yTޖ�;o3V�z�W�%�>6z�ݝ�`�ʆp��6���O��[!����f�����s���B�6U��^^.�*+�PF�D3X0`K @�%,5��������]���aq��}�D	���[�AL�3��jk��$�-2$�7�Ӏ?������2o{m�ր3�!��X`''��l��t�R΍g�S��v�ǚ9��2�RIc�Qq�`T��J�ȩJ�rEc��|DǞq����^E�xǧ�.��|�����jh���X^��|����#�q��)\�]�W�����f
��� �r��=��D�P�km������M��Q�C&&=P�|&2���73J�p��W�N�2 � H���#c��ֵ��9��É88E �)�-�RK����L���� �<���Xk�\ܛ�m�P1��K�HPR����R���n}|��>Os�����\<�` 5�C���8�6i���c�ͳ��ض�>#��BJ��
��5��C8s;M�,cE���(n>�7�H`<v���fS"d0�ç�
" ���	�q�0Xҡ�'�S
%��*Ζ�>n�\T$8�ٵ����u�;	�5A@����+_��4��|ȿ�rw�w�BX���6��Avˢ��T����{" ��<cX���f4%Gd���63M�k@�i�JZ����f P�\�:��ʸ��{N��ͭˢ�.������$�-���>�!ā��Pt�Qh`]����e5��8}��kٖ�1#�E��$���ӌ@�e�������Ǟ�;���2)+�����$2wn�6�T<�rD�˖�K��-+%�c5 pF�&�'��
tɶ q�#ѯ�l@i�n��mm�|*ݸ�#n;��
fd9�	�;��a�;�`��7�1�8[�3ݑ:p1���^{.$"��$u�-����>>=����+b�Ǚ�L󴓀-��ǒ�y��"@�:���%�{^̪�p�����,�<�SP�'�Qk,-�[����M���|�PscP���L��m�IKX�A�g�Ș�f�Y�`�$ݻ�-�k���σP��l��A�h����b��QNy���y���9��;�}2Ȇ��2�?|�l2��evB�-&�:E��;z�M�* �Xͭ+9soە�O������U�W? r ��D��S�=B��2�(����_~|�C}�c�C���A�rb�qp�ɲ0E�n3��@3VP��OE��<N u�v0a��j��ұcZc\j�36���%�z�q�����t�	g�f4���cGHW���ӥ���v8�[o�Ć�BΖ��:y*�8�X��/'�;>�[�]�=�6�S[��!����K��΁o�:@�!|�@�G=nr���yf���;f�8���l�n6{����M�[�0Qa�X��y�U8E�X��`e䰝��5Q�hf��	<��gl������� ��:pǸ�0�}�2z��;���]�a"Rp��'�j�����D0~�>ɩ��&�mn��@i�=�p&i-,�;�N!eځ&8��w�%�=������=�2;���(�o-k~{R�e�`�k鸛� ��c���Yzk6M�ˋ�:	����G���[�G?A�K�R��ƈ�����ѥ���| h��d<��PX7-�C�v���&�������y�%��ke�H����@�8з��;Y����
�t�ZP���	�$@� ���1$bf�"�5@( 	�"&���{�z`���%Ӣ��yz�����c߰ �y��9rf�.�>w�4�#_b��7(��b�  ����H��oQ4�c�r���ȑ�
T`@���Faz�0_��c�{
�g����!�^��<�d�ff�z�gϕ����z�ML�6"Ua�g��Hx�	3�U��>�>�s��f����w7�	 ) $ @!Yt^�(EB�� �@��D�),M��u�1Tk��&��[<��T�p갘�
��	�ù���U*���nr��tBXe���ZE�F`nR���ҋ������g&F	�˰8��څM�Ql�t��p�YeL"j�c�%(7:`��%R�ًh�D�&�6@���U�(預�K���mih�k�- �թI�LPsnH�6�൷@Չ��]-�]r�R�X�mŭ+)�t�����UEֵ�Į���Ml�5M_���'���tD��I6�2��5D �6-y��j�B� A�%��Li@ؤb	�%��!��V���^0��f��Ab��n��G�&�q|݃��q����
%�3y�[���3��2�v�/W�mm�xǬ��<��v!�-sǦ��	��M��tt Haly�0=Ʉ�C��y��-2p����>  $	�i�Z�Vٮ�}|��t$�I�?�f'U����}�X?�D"9em�/:��}ju&Kh�����e�-l���4m�і�Vt���k��<��Z�6��=M�����k0��Ps6]m���E���_\K��ɠ�c[�����
\%X�����ȄnV���c[�<�(��A|B�Xʾ�a<	"�];i�����G�XL	$1���b��.I)<����6�[�:��M�\�i2WyĆ�$�-GZ�"�8m̀�:o�:^~����F<P����|y������0�-��7�}_�W����	h^f�ۦ!V�f@:đE�䝧�<�4�2��� qXXX��׵�'�D0p�o{�KqƶZ�61�L��0h���~R�̕>�2�Vw�Y������9����>��j�P ������蛽�\�lh�vu]5�&I`�s�ɩ	�|X����	 �ͥz饩n�ʬUm�W.ll��+�(�=̬�����q��b�ǚ�y$�,������O%<�`j��H�x�W��<9 ޤ8�j;�"fe���,q��Q��y>��Ϟ��S�>���H
�������EfL�G�9��W�'�X�֢aoC�-`s*���
\������"�`�2UL��]�����޼�O���������Ƿ���#H�4��{S�e�I �Y�`�u�lXk ��S�p��-&7����d�Ɓ$w�]�6Uc���ػ�2me�(���GN�f����x�k kh[o�Ķ�V�Ka�c�OK��h:Ǽ�`A��Dc� a�z�	� >�F���N���������{��7"��aRxhwxz���A�&��Ӡ�$��	��\K.{P@֢���x2�i�6xw/=�a��Z��l��D@
P�ʬ��N\��_we�������|����fK����T@ �VH�>�<�]�7��5n+�L�uԕe����Z�g�u� <V�`�An�˭"�M���^5����v�Ѫ��o�&�Rw�I_�(�ج�k0d{�Y�b��ȑe�w,�6ڨ���h'��� z�-cB�v�P�d�dwpD&��-��հ�w�����q���=m?	a� L?VUq�ǧ��3�:,c���y�}q5�Yfv;��W��רY�- O���ߜI#K`�����ϵ�{��3ml����Py�O>tKa�.�{��ܛӐO+�G-(8'c�.��uS�&�C���o)���zD�#VU�#��^z����~�����Z��%���ջ�O����2�K�
8-�5����Wo0�eÓp��֤5��ΡO�Q��E�d���B�K8ˌ(D��U"�Y����V�?��o�2�y,O�U̜
1�'*�^��½W���:>V�aS�� g��6���wj�]@Dl�AcQ���Ib�WEhВSV5F�-:��j �CL'^A����z�?��0�U�i���'Jm"���_]�|>y���v�[�ّT��X(c,I���=����g�1Λ1aQ'���ȁLi���f��9lMDi�oN|DjB�k	ΓIlp�lb�&�ٜ�׈��2 �.� ��Ax�C�D�!P�N�,8l.�#��-��:6��Kq�z��Ę�cPh k����吢[H�kK�<l��@Hb2�XQ����w>����׿$��q�{�O��\ �x�X��f���i���%�fh�X���K�[�`����B:��6��L)&a��jZ۬�#4�s�u��� y�띧q���S�R�y���6�a�H���|"�i�^h��q��Ya >�A `!L�<!�I���pIDC�^c"8Y��$��n3�Ğ(�"��;�YO��p�Shz�-��K%�:{�`��B��zA��_A�b�l�E��t��6wa�upk)�D����w�/l��
̰���4�a�:�����h��a	�$ĬNoUM �����1~�5L���}U�	��7
a�z�I{���˶����l�5U�Eb�<��I�MM�-:y*�.l���lw�0�!�m���8�T���:����zNpmt��8���m��OW-)F��m����uk1s��ø�*���2��j�m�W=���4$i Y���n'��(�)8��2�@�4����D�z_�DD@-f(��o�q+/.�s|;묜���/�3�u�1J�b�#�\]R�e�GgY6��j��ݡb��\����m�'-+& ��ފ �c[R�6��n��[�����}����jy�0�@h�h�7�#HkM�'��3l[X���<	��%�����m��)�󓜉ye�-���"4'�\CQXc!`m��%���� 4Gf]������-�7O���#K9�̭�mpx��T� ����W�:[�S'��K�w�g��K23q�6��!� �;O1$Am�V{����;��
- �+��<��&(p"�0��G^�}�a��K��zq-c��<@��v���b��Zlϡ��!%�"��f�hSCsj��[�$�������$�F��o̡���H�	�i��4l��=��RÈ�@=��
,=��S�Vd[�|[4 `�EL^)x#�,�Ο>}������m��0@�e<D̼�n4�8?17��ｐ'�^A8�2����q-�Q�
b���O�I=+KI�&Ho�x�8Ԑ4���46>�������`j�cIQ��	T��s��XAkFJ�s�� @���sÿ�5W � ?f��s���8� � -F�59�s�ӷ��/�����/W�������7Fa�\w���=J"��B�'����S�К�R(�(I�.(��OY�,@��@.!=�y�LMy7w�8��oYJi\'���9FEP�\U�o��4U�Zǐ�����;�)���E�x�G��TM�E�O�o�qS�R9�6�7N�����?/�K�˺;�[�w�ڪŌ�"R��P���f[*aJj�B�EM]�AiKĹ#J�K��FP@j��DLFB��T̕��\)�ٌyv�hZ���"��7a�m�����n�n.�mE�Zg#���nH4�r����]�����^h5����M14��fR�XMIr<X���-phˠL��%��\@��e�%
�*�m�m�������f7\ �i�Mr�������&e��6ɩl���h[�Q�nU8]l%x;�=�+6a��+�U��g��2a��Z:��T����ۣ}L�v��vH�
(
Lf1Fj�61�d�וqj6��I�Z#Eqk�bۋu����Э�4�yyr���_�5 Ւ�R�I[��T"��
�3mVE��ܹ����E6&`�S8-�n�e�Ӱ,��l��YYx�n���6�wwtv��ٳ���T0�&¬�v�N}�X	#Ma�	�)~>zC�m4�m�"W�0�0lrY�{!��(-�j3w��K71�@`�4���h��D������E�Eo�rIu�w�'Ht��|h��ao�L �nn�x�Cg�E<��¡^�m8�8����Ζ�4�Y6�Q�1�c�e��瑥�� (�>pq��C:)?B0Y�l�2��y>����'�{���4m�@��egK�<t��<@�SPP.%C��[Y����`  �/DK0��Y��ּ ��r4�0��l��*��c[r���RN���+i�:e-�-���h���4��p'�$���q�������n2t�7%��5��K��d37���݄�L<E�ϿE�eX���F�qWkx]�[��5�i>ra{���b���hy���4l������>���mJA&X�oA ��2�� �d8�yow9L0� A���wrOz��>�Ͽ~{�;��7�>�$���EǊ+��e֍A�6]�W"FR�l��.�f�Ĕ�f��NCF��:�v��N��3���^s�<��8��]�����I���ró�r��{�������Kx�=�[������?����
 P��?eķ�e�b��0��~�w{�L���4����O-��`�p+ N�J��xX1N��QO�EN"Ë�v ��Á>-T����}���i-��.�,-!��+M	���>���ד(�euAޔK9Q.'���u��D����[���if�C�rǳ<@�n
�p��:��tA�����h�wn �c�&���C��'"����u Hr����{�>�|�9y^4֮�`ꤕ(8S"t,Xk`@`��ܲ԰���^�$'n����N��BI�E^������z��i���ԡ6�x� �e�|�����+۴ ʱG(����<�<�����/�d����W��C#�i��6�$��i�r�����玖�4�`v��vi��e�.������ڒ$�  �6<D%�AD���e�wwS�\��Ӷ�*���U�A2��D	BW#0�h3p��&1P��,���c���׺�,�&*ȋy6Q�Uj9��M펜�T�����r��:�ޤ���̇����ķ�F�Sn��4�s G�1}��d\�q�ZZ�\���r��w���m�]qnUn�����Z@��4@��ˁ<hn������2�]�HrUx�ˇ��K��`<��M�8�m0��WSȐ<n�^b1^��{o�.�z��@PF�l��W�d���Q!�Ϙ����~zm,����a�)��j�x�U
�9YV���WD��1U/���V�UO��5sc���:4|�+�x�r&�;�e@1RiNg�ڢ\�b�;>�{ٵ��j-ըyQ@�����<���mX7:��-e���E�7Y<��Q�fnc <��yx��%����F/��IP��JQ�(�x��Xw�F�ox*�(�V*�1LE�����cBFCIb�X�m��H&��F�*P�cfL�1�#�k !���� ��3� X�mC�, ��@��\	�n�t�}^}�~��@����*�VC�bRQ@<�<i�����m�N�Ί�>�ۉ��y
(m�-|��Z����af C�`����C�A���Z�,+zpEb�j�ЊQ�IÄ�D\�/3,��S���7���;Y��޾�3�4��L4�x]��i>.ԛ@��󼓦�����O��$
IDH!g��&@��F��/>3x�D����L���L��À\�ˠ0G@�2V��i�ѭ)(�B3M-�顈�ʪ�s6[]H��]͕�̝>-�T�Or'�0,�X���눉�U��l>�Q"ǂ��]� @��';��\�U����^b�RMݻ�P�9x&ӗw�wi�H�2� o*�	�C����z����]f�Ɋ�]��|}������L�P ��s���P[��d��Î�Z���m�fdAH��m�l����,�I/���z�a�Tt�`\{���1jcC������Ϲ�b&�T�{�=��ahpO%�'[U�b��r��X�Dy��^�p��	���"d2�#�c�2�O<�o����2�j�c�hN8�~ŀ��>m5� �|ŬX�{�����"d���h�s�f� �� )��c�L��2���;,����� X��p<o���-�IoBmk���,P�;��$��X�� �Os��ݜ��S*w{}_o~n�p6%����	
#^�a��LM,��^�u˕��4
� �U�.ej۰�L�Zj����+��l9�(B�8�F� F[��tiS:]-��M��Tإ�4F�묟=�!�=��z�|�{��MrE��T�^�����j`,��e.�5��Yڊ���?	��9<��}ᯘ�~z��UF���9F� #!���`Lw� ��U{��[o ���*�k��qŋ����	A��o�����:�Z���U7&d���6��Z�y"@w�|���#Gs��;ѡ50��h8!v��+Jb�@uLX>�֟��!0&��<֦R����v��酛~5`�g@�:y ]���j��Kl#�ũ.��e�~Nt�T<$C��!��LȀ�J2�7ki�)����z������x����^vM�0�	э�x,*��"�l�x�+�L��L��T���"I1%��Yu�s�yqNF�<��<ɗ���-r�~��4
��xu����8x��P�f��a���  �-UŁ�>gTX>|��E��O	��2�9*e�.@��xoe�����f�~��V�V�"�R�6��X֬f."-d5k"j�B#	��b\ơ��[>��3���sK� @y���jϱ��-�\���y�e��R�*�[Ǘ���yK����^�p�AF^�(��'=�/q�б�n.����\HŞS�k�y?�9�iz|�&�:U7V�${��}q/rc)T��� �d�P��y�KDe���)��,xR��c��NJ���٫�F�z��^��+1F�TIb�U�1,��DPb!�\ 
��ֵX-!� $Q0�v��\0��@"��b� e�(���ݽ��MW�)��يhƲ� �)Um%�jGde�̚��%a��M��K-.�l��VR�]��u3�֍\�T�]tu*��B`���j��4�5�N����Л:	�
P�4�M[1��"�K\;���e�s�܌rfٛ�΋�е�iZ�nUk3��B�mca�њL���X;X�Z��vz�k�&������Y(�]lB%�4͆�n4��V�Ms=wτ�$��@1 �Ld&����8鯒�K�`��M̹����1)�DId�wш��&J�f8f��P�kRV�����S�Nk(fХ=a����0����p��j�Xn�]>��~��O|��z���h:l����­.m� Sr6����ja$i�i�L�~y�6������;�����^a�	��/6"8%��;
�X�): �>�ۉ�	$ѻ08.>̂T�`�$	"9;^g8�i!Z��6�0W[�V9٫���aN�@�pS--Dswe8-0g�<Uveb� a��w���_�~r�-�l�	�>�kga�n}ݿ)f��iq��7K�*��w8�a:��M1nc����<���R�͵â�EȌ�d�ܪ��t���>y�zc�w\DKx�>-g�<�}qM�lel@�:睥_���,���f�$D�q�{�3 �6�VT��E�)"؆]��l�U�ˣ�[��le�ʻ	��@�V|#y��c):Y���[�<��a~B��0U�� 4�q����=l����ޫ;��=�=� ��B" @��1�i �=8%�����O���䝂���dn�&SZ�h���h15��Dvع��l���12�]�o[^m�T��m�G�NNL�/"��[t\�@�O���<��z��'�-��S��50�T2oA[�xѲ�l��]F@h ��I�;WZ��}n�@;;�1�(Ъ����&��S�x�c��h&W�Οn;V@�k�4*�Yu�(����fpdss��E`�1��5t�,�h:a��'H�sΗ!����p�c2�"J!���a�$�F"�KA�Yo�~yk0[Ƙ˷�yڀ�0i����8wn�*���!i݀��$�WN'��RogC��7 c����N��
�8t��'��ఀ���5�;��m�3kK!����<��t�b�Z���ʀ!���'���&D`K�{�*e��ez�?[��Ҹ�e��Q�e�Ӣ�Z�̻6��y~_\�|㼼?%�|9Klc������3���m����Ki|@���*v[Ź�]�� ;=wK ���ܽ�6K�w��xߝ}�:}�~|���D���x��҉n�V�ۘJp���fb7d��b F6 h�,Hq
=���	�N�]�y�V<m�BdL�v�p�y�\��Gr�y�5!��gm��i��h6���a.Ǜb�d� ֒awC�<��w?,��}��Ǘ�|Ǟx��qEJb%���[qq0���[��cG$'�漵��]�]O/\}�0f�� 2w<K�d\��c�Y��zy�~�;!B[[��Μ��Eo7`B!��w� �id����w����������0�z�����`�oK��zՀ�$���:��l�x.8�^z2,����7������Av=y�aS�٨ǫU>��^vyO/a��\�fLЙ��xV'̗�ʇ%g�ꗙ9EJ�LԺ�(�{�xz�ϗ��ܿ�z��2�&�	��1�t��ޕ�-Ue>yO~��~��T��S�[ȹO с~�����Sֿ��C}jm\ߜa�ʝ�]� �k!�b@N���T^Aq�z���&^�����qn���E3-�v�����y�<�<��j��Z�0�5�����+ y���O���@�[v��t����G�/?<�S�4���nk|}X��u�
��ڠ�^�8@�;)����[*�*�&F	T���t�l"Jl�k�-�O
v���A�z3�
:E����Hl���0CE��5|�9��ϲ^I��|����3BH���	?s8$�>7�5�_]��8q @� /7#K����ɛ�:�&l��ښ�ȵך�&�b�j0*��6���!��o6Q��\��k�.pwx���1�9Y}j��,<eә-�5O<�`[�̨��1���BΜ�@Y�$�q�'f��;�t"���"E4��.���/��,/�nz���eā�v�ƸKk|��^\�ꑬ����ػ,<�u������# x���-$i�,7�[p�:YsS��;��A���f��dͱkݱ��Om~\�u߻N�N�pz,<Z��0Vs�o���|�;�]d�%�n�<��>ll����ӌh�j#�;F2p�D�.�"�R��]��k��޸�#��I����3����7!P,2��H=<�gM����C�܀Lt��ب� ch�c3J���,�c��< � `3���U0̎Ev@ZKv���>l{>m=W�6|k �WO!-����YF�*yM�P@���`7��'Kd�O/��󧞤@!!.�&��'��G%)����DR�P
���Z��hne��2��L�u)����tnX���H
���	<�P%�*�5���7^�J�+M�Xx������[�0.ٽ��́I���]ň���O-m�(������aeE���[��p偞!�R�f\w.��l�<m`A�0�nw�{��X�i@Y���
|��ˆ��[������>�3��<@�k�Ya'Ƌ��)e�m �o{��p32�Clv���%f�,ҹO9��~^�a����(�ͬp[k�$"����3�ħq=q"�2�r�zKaq&����d|Ǽq���Oi������0�wE�˻ޫ��¸�3��O>Y$��T�v��x�cD6`n2�c�0t�`�	��R[���j}��㻝7j-�ԷY���N$0��[H{���/�V癘*���	n��Xx!��� 6�%߲a����0h�~S�@�6ܚ�h��69Ya�4�~�e� X�^c%�ƻ�D�C�
 �"��Kܑ,����P"ƀ.�cT�cB�b~�8�"
@Ր(hĲ�N���N�7'�����\���}U�N0�bɷ��b"&�u%�L�SO�!As0�������L��p���W�zT�O����c�'j����I�20���,u��Q>>w�{N�#,d�sg��b|���D׽�S�eS�=�c��z�q6aM�A�0��J��.�d]��i^��^=�&v�<K�'e��u3����r��9؀��5`EH���m�E@B� "ha�jX���7��X�� =M3{�Z�+(���X���q��M������`�v]�\1��#4�V$�Ѓh	G����bK�b�jhX�қ(�-�il׫`���Z�Ţ&��P��.s�f�����&
].�M@m���ҝ��[����6��l1v�ict���Y`��)4m5�QA�;X�űԛfX�`��R��0h��Yl͙�ԫP+�l�sb8�i��f7kܦGgfjK�c;X��x��0$@�R�E��ȉ�빢H	��q��BI��/��6�M$�����䜗�D*Jv��ؓ[w��ن�l�mŭn��P��Ѕ��X� s��oRVR�Z�R%��3-�ᷤ*���x��D7��}�|R�q��^a֫���6a���w���Bπ-r	�֟���ׂ_N*�h����X��p�e̸]��X[1�:۷�Ӥ�D$�$sf!�&�}��G��9�o� EÍx�����s:a�o�{q<nSx�>��Dsc��h[�e� �]�($�v��4[KQ��W8�=%5"1�D/lt0�QŖ:y�s��p�U<�>�#�O>���`����v)�8�˓�/���_g��������h9080-�T$K� I�-÷����
������]*[L��k��\	=<�0�0�y;�؉��b�U����6���t�v��~���,�5��l;�'�b�������r� 8J��Yo�y�����@N� ��i��, ��ط�
�4�ri i�^h��y�4-,�y��T�cF
���]ߜ�zyw~�|��3�w��_%|�PR5Ua�V1t�QR�a���ptي-�u�@�^�f�9G<�M,���i2ڢ;�d;�f6�Ǜ�8c,0��Z�Rǈ�a��k(���]n0Si�Y3�%�l�+_�	�P�/#��~�Ш�>�onr��Xgv��01��T�ACk,�Z�>����=��v_��=� ���||(��O���j"�v�z��]k����'za�t޶�<�4Z����s���؂y�bF"O"`�"�����`��[���7%�F�*�j�R��x4��a8�c�;f�'�m�;Kd*�������	>���#|���6���ij���I�D;�p@�&
�q�r��ٽD�އ�0�cUp��z6���[����X3�6i�r�u�:ky����<#;v�gx�ZAv�ٚ��PO�������K�c
h�+dB�YZ)��7����m��f����ioB�ʓ�����
 � Rdm�~33_:�^�YFb'K��ʿY�z"!�0"""
����\8�(.����GeΌ�#�b[ad(f�E!��U�:ݛ�Mu6�k*�0V�QbRI�w=}���6���������;�u�V�42O~vo+ �f�WϹ�[m��}�9͎�;bV�9��\6+���������^w=�����1>��dW��s���o>8�a�HN��<�8���W ��ZDȃ1ƃ]m^Yl��z���=��d�z�uv>���Y��ܫĊٮ���(�ǌ.�3Գ<g����	B�����M^��N�w��}�Q�*�SC�j�[�{=��2�d�>ۘ���E��DY��U!6<�OI�����O^x�>�xx�ɫxl���B(�\O��H������נI��QYL���\S��`��Q򈢫^�ʪ=���4�
�v�j�D����M:S�I�TJ�"��bA$A�OB,>�:@%`$�=E����rM2)�CL�4�L@�F�s�I1�e%$F�fJd̚i��4�d��)����2�JY�M8��k4٦f��Vi��L�9��)�l�2Y�M�nie2�L�eM)4�6K%s�q���M�s6"-2)������b���޺t��9'o4	-u�����&�}��l�f ��,�C3+s�{껯���T3�W�n x�;�^շ���OZ~Ua���\��A��w^̲.NlJ<�����i��� {�}���b1�N&T:uqp�R�(͹�$���I��/R�y�/SC��\��|�`x-��Ctߡ�Z���S�lv<0Ձ Ϳ�vno2g7{������ߝ���%�s�|����R�*0���0A�mLK���st݆1 :̎�,H@8�ͷ+�J]�7M�i�F%*94�K/.F����|�d��'���l`-�2�N��96 w�4{g��sP4y���,0�Lf���r���Zb놡+3���,k`O�OV<�`�s�Iy'"�jñ:�Uy���VJ�dxL�� ��U�X kX���b�m�D0k���ӌϭ����Y>ܹ+3y�K��,/3b"��&���G�����Jm ix�W����
�^��^
�[���2+��U~���a��0�3 uu��+�_=��{*U󓜩v3,�K�6�IED9;ی�vH`N�z-�`I�D�}ێ���d��C���p�@�a�ax���[`�{���"�eS���Us�}��^��y�q��f����C(����i��s��f��dX�zWCPo5���5�
�7�\0�=u`
��^�K��1	�d]l��h�	��2�L2�&gϕv^K��x���T�B�j"�i�WaD�UK^Z�֥�f8H�K��a�ڄ�����6"8�9�#+O��d�:�fN`�,I2�*y��өO>�3�
�9 xw���C��Z������
d���nkm-o���[ ffXB�"3A�Tn���'��ԓ���;zktQH��W"��xt"M�6w��ꗎ͆徸��Dn���X�9���zx�]p�`	�d�p�p T�H��J��l#t�;�#9>I�ϓ�Uˬ0�S���;�CO	na�^�E�9׷^��=��ɰbߟ���W���VÛXX��b,2�e��S�`x�T:�<Dz}mDR�>�{���L촞4���A�X7m����	��� ���"�+\�'{7~�:��ӑn��s���>z~���w����Ai��.E%����a�L.�p9�4K�p}�� �Dn����Sy�
�!��{��v����>q>��"L4a��?���,��k��� k��a��I a>�~���L��Cr`i�`g���@߀j�����������A��EK���i�f���.͙�>�o<��)�$���2@&��i!6i2$�7��!�d$��0a FB� ތ�#0����M���2HU���&�qm\��&��	���0a ��3Mm�FI!') �I4:�$	� @�@�$����� �@��	�I!1@1��$��L�CLao2Ii! �� YlӒB#	�l�;&1fk掦����2K� t����ׇnu wC�u������C	��r�j��%y!]π�Z��+kmF�mm��A� c	�ՙ	��#�S�q��v��:����gy:OV��Hj`��'�K���5��gp!��hg���`	ǜ5vv5���ć�&���&�����3���0��v{ṵ��,P�������/c��8��y��?��9߄;C�gםO9	 ��z�?t�C�9'C���q�����` '��"��@����&�c$��}��u��C����n����$�zϐ�	�|��	! ��5��d�I�됇�߉!�đ�=�M�� ������?���~�U�xU���ؼMy����+�Wj�(���p���}=P�ï_�Ԅ��xHRtrOc��:d�V,�!�bMC�����ɒd�����5'�'��D���=�zt��q�~�<�0'�|U�d�tu�����||`��0�Mq!gꌐ�N�P��f�( ʯ��(6��w�C4fa7�}l)!Ȩ��ʵ�el��Umɩm����skt(�U���%k\鳛[[�[��TV�-�X��m���f��,�MSScjk6mZ�cV��ũV��kUf�ʣj5lm��h�5e�j�l�kM�kVl�jl�Yem�+l���e�d�6R�5M����\�3i�66�TV�Z��J�*�cU�+i$��! )�		�Iǯ��`ŀȄ�\�odL㱇H!��0�7�_��L�u��;�u{0�C�����b��������C�H	d��@`M:>s��zy~Hg�������+�I��2u!�!��I�HJI��|!�ɯQ�=�2��>�R,�@�7����a�O\�=�{�0`��C���������g����B}�z��8}$���?��=Rh�q�^�jm�vZ-��,h��E��4h��ō4i�Ѣƍ�64�1�E�4X��Dh�bŊ�4X��*,Tllh��Dh���Y4Z,�Ѣ,Y�Y�f�4h�,h�h�cF��F�4h��F#cb��cF�4Jh�cE�L�ѦF�)cFƍ5K4F��ƙcQ�ƍ$�Zi,h��E�#F͛R��E�4�4X��i�,�&��Y,i64h��Dh�fh��4XѦF�4Y4X�Y4Di��X�X�4XѢ�e��ƍ��#Fō4Xѱ�4X��cF�,X�h�cE�E�ѢƋ,XѦF�4TZ4XѢ4h�ll�M4hƍ%F�4�4lF���4�SF�F�2I�M4X�bƓDY��Ƌ4YM�Xر�bƋ4dѱ��ƍ64�hѱ��Jh��,LѢƍ�6,X�h�bō�4Y#F�,lh�,X���d��hѢɢɣE�)d�d�Rh�cF�f�E�4X��h�e�4X�X�F�,͋E�F�4h�X��X�h�E�E�,h�F�%�%�64h�ch�SFѴ�,h�3E�%�%�ɣF4lX�cE��I�"��E�%��ō#F�,h��,F���4Th�cF�4X�d�b�F�,h��ƍ6,F�4�4li4FƒƋ,Y�4I�E�cdѢ�F�KK,h�X��4h�bɱ�ɢ�F��Œƍ6M��řcE��#fX��ccE�F�4�,i,Y4XѢ,i�,h�cI�M4�4lX�b4�,h�b�bɢ,h�M&Ƌ%�#F��œh�cE�IX��4X�fX�bH����ccE�&�,X�b�h�b�4Y4Ti&1��B%,�&	1�F��"QE�b�ڋ4���9�����d�t�a�'�	̐�	4�h�P:l���=$���gC�����	��{�SGC��hC����!�l<�_PH~�φ��ϢD�ROC�?,�|�$����<;I�A>rFC�9���1S�|d�Y'�����C����=K�ß�'R|o��		$�x�� �Ha�L�C�C��H�G�t<O��/��Ԇ�gB��'?��C�'��?���9��C�f@�&:'B�!�{���D&S�O��C3$��A`��|�)���"x|Hxy�?���&�s~ {  ��D�����~|����,D�8q���l���~È{$��B@�!�a�z�I $� }�)R�d�rD�����|>b�/�ԀjCRx��a5&j�\d�sP�@�#�L�@��g�۶�u��:�!� ���$f�Ԟ]z��Р'Hj�Hxu�מ��R9&͓�0�O���10!�I�HI$� M�gs����0Hzt;}?q��?��q�I ��c�!�I�đ�d�}����	�O��C�v�:<C���'�f�?��C���9����t{g=��&᱌=�I�Ol?9�{�Oq�0�����>�'X|�a吟��!�%ޡ �B@����������<�B��a�&I �7�3���O =x(�s����i��H0��n�� BBC$��m�@<�u�!���^���9�<~b�����(xu��	����JB��#�F3Z��e�>0���t����b����0�T�����2z�:C��"?��ݮ��go9����̈́=g=��C�%|�A��:��0�d|:�:!������K�86O?���I	$�d��<��&��s<͇��=�{љft�WP�:�B�c��&B�9��h�2O|4M�Hj���xD~��'�~���5'xN�|A��,D��{fa�S`v0���Xd<���x��֢3��Ï���I�|�����P'��?��L�o�d�I O�J`���� �7!�G	'����~��s'�O���S�$�@���'����v!�a���N�>h|Ф��	�О����'#�ua�C������h�߇���i�~��}Y����=��)�`�5Yu*�������.�p�!U)�4