BZh91AY&SY�([8	_߀ryg����������`�         �          ��$�@T�)AD�8�E�R��%�����T�����(�9۝Q�n8>� kC����
:N{�(�G�o*�;�.4:(i�������>>����h����E��|\���>�}f���
>��Oq� >��=�c��M]��
! ��:L���]�(�Lw8��.�O7N@)3� 4S���#aƎ�9�(�qf��/|��>��E
��th��.�Z�$��           P I[` i�)R5OR �h     ��T�ʪ��0�!���1i�`��UJ��        )�TPҥ	���h�#	�&�a����B� !�d�1�4���4h<PmA&�ڢ)�jd�!� � �:G��{;^�����s��I�XG{P:���
�@sUUz�D=h������5DK�D0?��������o���4�:q����dcm���������]�p2����9�sw��\59K��?�rG�T���z��]�r`PUP?<�q��UG��S�Wϣ����a���(	�_�^��D�`��L����#0yɪ��/��P� �φO�'�=�ʆaw�ΐ�H ��L lx����}��Lo9�}�_'�ɞ���5��9��k�Gx�}{������ߦy��[p*�B�PPX(%�����j��`�B�PP��
"���B���1���A�*
�
B���p+
�`��mЬ-�B܅��P�8�/-Ь*�v�aPPV�[�XT����V


���PX((,m���PPX6�+
�AaP�n����XT���q���m�v��
�AT

E
�`���!m����-�
¡P�(V�����Vq
\T-���T
��(,-�B�m�AB��T8�B���

�
��
�B�Ơ���q�B��+��+^!�[hV
¡P�*3*m���
¡m�[y
�C����*%B�XT-�
��B�XT+p*�T9�r��m�T�T+
[m
�B�X(V
�aP�q�T
.B�nШ,*PPX*�I_�ΐ�Ht��((%�T

�j������
�aP�6�aP�q��
�A�*

�m�+
�aPPX(%�m�wwwwwwwv���X(T�B�XT*��賡�Htä:B����W�(¡m�*

!XkP�+
��
�p*J��!ơP�p+
0�,*�5
�`��Y)p*rqp+�aPnanC2ۻ��P�5��XT*�B��q��aP�y
��¡P��(,
�9��(-B�XT*E
¡D8�* ����۴+
�AT*
�0�[�X(V�m��+
�`����Ty�b
�B��*���0-���aP��Im�w�A�Y�u�CB�XT+
!n`�Pn([x��¡D*��R�-��(c
�aXR�V
�5
�a��B���n5
¡�J����A��8�[�X,+==u��hv��!�0�+
�B�K�X-B�XT(¡P�
�B�p*
�aP��D*P�V�*E
�T*D*�B��T+�T*�P�(�aF
¡Xk^!�/�XV
�aF
�Q
��
 ��!PD5�x��B��!P�*�1
¡XQ
�aP�q��#
�aP�V
0ơP�5
 ���Q�T+
�aD(�aD*���:�wv¡R([�XT(��*	rB��ۻB�X([���wv��aP�
�T+x�`T5���
\
�`�P�9wˁX(V�
���
�wy�T
"�c%IR)q��  |�˒��9r.�~k������x���s��?��z~��E�����_��Iߛ��fI����0u��<������3�>���@~��6�`���"L߭�H����2L�����?1�T�y��\�(�X���ԜqoN�W5�ꅣA����&�)�9����uJ'Ӈ�#Z&h����xW"�͋�E8�gd�(�w���`���8(b	H�6X��R'&���͛S�O
*y.e��;�w���� C�܂2�Sʋ^J���&k.}4#χĩQ�z�2]Dٛ�B�Nlw��"���ˠ`Q4o���F\�U����1��T)���b�|���@�/�uQ �dd��5p��1�U�+7 �()�WV^NM�:�A�D�j�G*V*��d�zR��<P�X�$M�P�7p��Yq>�{v���e�ҥQx⤟t�xz&��f���g^E8x��P%E����Zz�b^T:̜��y�1���19D\fP�Xf���-2{{{5D�c���.�`�!�9ʷ2ȼɺ�w�4�	��Bj���!
q����g!ėx���Wr�P�"�xJ\�L�,��n�DD���h����Ũ��5�^=;��ʅ/O3� ��V�<�Qwi��̉Ǆ�N��3s8e)z�@ٷ&�/g
y�u�Y������ȸ)N@���P��4�����^]^%w%�Ҋx|R�M1��b^0F������B��9Hz!\Z�2
�7��B�Ox�T2��-�1��2���h+F�r��U��E=�Ù�䂐�1"C�|"(�<�wr!��TTE���{��*E���e�0�$]Q˦�9X��Y�V�|�8�Y��B��3��Lj!�FbC
��@��E@�ydb��ӑ�8%
�I;�|V��u1�r�̧��&��F[�.��J�Ž�T�R4�(Q�e����!�lP�/�к���sOB�3�&�Y-*R�
x��{�9hR�"�;�8��o�bԌ.e��T*���X�'QMo2��Ӛ�03 �!A�R���!�
����vʚ�Aҩ2#p8"_"�;)3����WOS/0� ��q7oIA&�1S��/%Dd�n�e^Xd�2�TxŻ����1Q�Q0\{/&�'(��E�T
�-q/u3�T'�s �(X�𼩼��ȷuP^�\Ź|7P�
R�DUɲ^`{�aȫ�'".�݋/U��P9���0*rj_ =U)�Wx"p���".2�<���EQp𪬅W/`���U��O&�(UF^�w8&E(r�J�3�O��|���0#x�0C�(�w�Md����LľN^+�w3�^f�˱r��2��UNrhQ�V��7��WRb�͈572��U
�è����c����I���zyP�d�F=ы�U��ͅ7�4nP&�}k.e�#��]%1�&���(e�L>FD�$b�Xz�g#�HQy�����(T�I&��"r �Te^+�5�(��%��f\�D�dJg��fL˹9���&�I�Ȉ{&EX��6�T���0^��]�B��$"�'+.bB�.ɼ��sY�e��SjL�=��h�̺)�&�B�B���O&���z�k,���b�C�ޞZp\ӧ�@������2+]P������n�3X*���O8�fi�#!7�lbUJ������R��30>_|�'��{�0�i?��wM�77stJ�  �`� S.�6e��&J	v��  �+u� V��	rX �HU܀
�7@�` �X*  �%�J�@eeLA��
�.�p))  $D���b�Xبa�D�ܕ6�PKD7wkD$Z`K�Y4@� "�]���
I X�Ar�������
a[��	���ӐB@A@M�dF�E���D����������f��ww B �*�D\��a����d����Y��ϝ��[��]�K��b��,���]��>���1|��������Y�c��9q���p��{���z5�N��+��:N�����\b�뺶3���c��G��{'�5�ҕ~]�6�S��J~[�Xm�bx���������=���wk%�"�J�3�v���cg�����iü��7P�c�9,(�z�<���T=l����淠6]=E's#<��@�an�+R�+e�鴊3��7;�ݼpm=uqt�e�J�]��o�޷�]���$6�	��I��bFԞc)��s�=1��	N�k��^�b��>b\�K�ӻA	vKm���8cn�:ޔ�FsH�jy�/9����5�OX���E���3��&�3�#6���Q3��X�Mؖض�`�>;�Dlg������U����S��!�z�5�nG�!e��"j�6�Kg �(��/X��ԡ:�\�z{<:���˗��r�Hղn9�Ѭv�fM���s6T�=��Ɨ�^g�ӌ��l_H]kM�gm��]n�1t�iq�n��=l�P�z.�<v��`�L��7l_�;�ϝ��n��buE��:|1�ݞ�z5�s�8#m��<����9]��v勄a-��=FG<�eLqٕn��!N�^�U�k�텼]�:��$/G���ڰ幧(�9���w%��rs��ө��f`�@+��g���|��]�\Z�lM��]E\r��H]�vy�V�d�7tV�JBh�J�e���0�X���n�id�����7�|<��qv-m��n�B��\.��h�h2A$�*[��Epr;'�"��+r���%Z��qt�d��=�H������l����b.�!�D������z�[�X�b���Z哴?�<�Y�*L�X0w4v�+�M!�be�lFZ8���*˳j�}a�#��n���o �и�]Lr�˯a�e9�3#ԑ�u��g��y{vz�t��k�]��%zKWh..v;���������+�V����(6�c���e�%�Xۈ,��V�n$1�t�ݷ\g��y��%��3��A净D*�r����6��r\v���oOf}�OF�`�/^�'N�r��/r��y�p`��fM!c�$+[�f�G�˩����hzy�*q��K�Վz��]&�c-��i�x��#��v�D��m�.o��V���6H�k�t˚#	�mHntJF�d*8P�(t�?�߄O��~��$��~���-�?� �{��������\���"��nw�5�����ય����AͿ�0|���<���p�'+�^�����F�.\����w���8���?FM��d�3 ���I��5�oy�B/9����
2�E�q�fk]��9�ZB�*a�.q��8���4��#䷔=��̏��Y9x��I<���Q�'�#����H����Q|Mx����=��_iYh#ǩ$���CĂ�f���8�y��x�"���V0,"zBOgE<��Շ�<�#�N^ӏi԰�E9��Y�l�o<�p�4�Y��/#�B�y���������<}$||�����"�T�XUH)�^.��A2L�`H���
�;Ǣ�_�[����|N�M1x����D��a�B
�m^7�hET���(O$��H���v�2߿'R3�}o4��g���ޗ���������6]ҧ�4ha���Q��1!&���0��.� D�(�T��y��&�ZJɧ3����H�-����C�z�`��ȱx�{x�-�e��B�
u
��a	�����d2�L�5�3!E��$"�9���P>L��3.���@(�8���"��_{�o����5��,����>���*b��2�ēp�<L���1�%�8�!���ªE[ς2�=�L�&$㬁X�<gt�`��d��A�hp�&-�޾=���
ǼMOn{w�	�ѓ��l�2�]�V2Na��}�OP�P����G���� ���{��rs\[dz����O�%Ϣ|�F.r��)�K��ȇ�w��y�&�%iRH��O`�����}����?���g2�W��V?�IR&\�()̋
&-)!�#F��^�A.�H�0�Q/I܄Eʔ�|�}�ڋ�E%ksO�.#�!�����OH�j\=C�Bp}/AǓ��LQ��u�6Ie�+�4�����?_W��'�K�e��~c>Z:i�~��Ҭ�����B�ʞ��[;�|ƿw����^��y%�!��{�*O`0���S�j>�����{�oT� �{x�o��f�<��9����#���bL��2�C#"U���q ya�08$�K�by�L9�-�b�$�r�2pY:</�#>�R�@�&���}�~'Dw�w��V�s!��4��s?P�=F{�8�z�}9�zȗR�q��3���C]B�����Y�%C;2
�0�ÌsB�M;�C8���c���y���x�x�*�@H�J�]�%s�Y�>�t!=��c�����+�nɻ7wt7Y�� ˢh5d�	!��%h�!�AX`�#vn��@ 5h�dPM�Tj�m��x�re��߫P�����������}�	�H
��,j j��W(�T@P
YM&�� lٲ�� .����(hi�vn�Ry��;�Y/���ߞ�Hm�GS:73���� ٴ<vY�7��u�=?%e���bݫj]�e��u�q�V x!0"�m���[�9�� �rX��kz�{��Qj����h�-+��E�	ж�
�os�ֲX �[=ڒ��$t�\�oU�f�.n��k����6�Y*WT�7�U���%���\����S�a��cc�W�g���ŵ9̛a�u�tYy����msũܶ�0=�n�ܠl����|����;`v�AH�H�(�+B% P��ċ��uNW�ȱ^��MFe�\�~2�ٲs����/j�w��VE+vl�3=ɜ^佭��0SWJ���a36�o8�/y0L=f���m̮)�9�GKp7�d�ml�E�c���Ii�Y�ǐ����C�X��8rQp��	����~XoC��uO����ͱVg�,�'�>�Lޯ8lk�)��m�pZ[�a�odŀe�T�N�٩m։*�3Y���}��Oܓ릎OQ�|h�	ϊ��Pf@�`����	�i�x7na� �j��L�[ki�-�>�
� �2�"
�Q	<B�x�CT:�}}����T��X�N�^�kݍ�>�N,����W�CM����bk<@0V㍶a;>��D�b���k�E�n��z���Rg��Z�xz���j�� �=Z�����|�^��lQą��Fy�˲o\*-1�Cu�[��6�hl��y���2M����u�럛���1wiz��@���w^�=4����1@z���k�Z�[�b�>�$
"�f?yW�˷<ɼ�̝?y�\��g_��w׵��������O ]m6�b�y�s�ao	/C�/;�v������V��-�,�ŧ]�B(^Kj3S7[�����~߼�ԝ�]p��m�o۸}Tަ-�vja�?��wIVۍ�O�����pIE��U-����������{��`Ic�v���{�wH�`\ă�{���F�6N��nߜ��yO@my�L�څ�io4��1`yB��|�&��^�����u\O.���~�Y�|�l/KT� ��	|x�]��-.�h��kDd�k?�v��t��_���W�Ug9��k�ja1�f���������S7�5���a�l�}=3z���u���DN��,���<,��F2f�] e��n�f�V�@[������3Z�uɹ�*{�����V�ՏGm�i�M�V�oKXVh%�kʦ^p��ϫ�,	oY���FD�&Rf{�۟]��ܻ�ߎ_w�=��]M�S�*y���rF���Uu�WW��v��lj�t۴�%Cf6��<���j�T�2$Z�^ e	��f�G��v�8�b��6��e�" �� ?O�h-[������f�`H�g!�K_F�3m�O��Sz[��-��=[Q�^����-a���
�Q�<Ar��*�z|���'M>�0�P|\�K�eu>�Y��_���uQQ^��5�
!��� A@#���]wι�C�QoO�ڀݝ�a-��@�[h�[D�����<Ct�LU�O,�;$Æ��4��{q��=.̛��p5��$����rq_�V���I�,��y�?��o�y���3+�$�=�fL��m܊���$V>	w�Ly��J��]W�z|"��ا�)._�y�&��L�Ņ�Ag�Ib>G�5љ�yx���ʿF`�x)�'/oرO�4J&��_}���}D߁iu�2bc���c)z�s4��?��z�4�(pD0���"�U پ���@@����X��ŐH`KE"����uc��7�����$��$��\��c�X��x���3�����X�h]3�׽W�zHӁ��ὗ<�Xc��?�䯄� M�Zh�6��3lŀ`�i�-���������lc�����&���"���7|Ϥ0;q��3)�2���.4�e��.ǿ�z��c�*�~�0�[J¬�l3����BC� m�Y�[87\�T� ٝ-\�w��׷_�w�}����z� �%�"""!C�r�ꍠ�e�F�E������)JMZ�oY�0N�����iv�p�9d�b�!d2+�)%�,���㐷N���?���-�R[qv]�Bɵ�^��3߿}<#�Hq�eK5��{��O fS[jÇ� ���l�8�Qk}�N�|-8��Zp��7����ʄ��/��O����f	L����m�y���	�-�AZVK��j �$��M�O���l@�fG�_�����:�N��\�2;���U�s@>Lυs�u�7GSZ.V]=���~s��1~f�""t�cd9�4�\HE:��GP�H���/�Ѓ���oz�2�-Ly�d�;I8��|l�y)�>b ���������%��n�n��e�΃� 3� ʚ�a?|���Yanh��GHm�m������n�`��m�HZ�5(;8�FD���5�I� 0�M��v�D4� q�"F�k>�����wR_7�ȼ̄F����Ĉx�j��-G�apw��e��`el~� �e����:ZM�t�!�v�B��T���Z6Vr�<C`��}�L�"\��A� ��w>꧳��oL�ϻ�e��y�]ԯ;ﰺ�#3���'�na"G�!73AXjB�=��!���5�E.1#�Ӛr:�ٖ��q���c,vCjV,nǇ�i�c��I83_}
[�����+�M�����[��c���bC^�gKCb�<�t�[ ��m��R9���L'�ٍv�e�Zn���{ߍO�}���#m��Ha�q�<@�G=nr���yf�a��gl��xD[ ���`��`�L�Xm2����c�N����o�������x�5#���2�çxqL8�#������� ��:pǸ�0�}�2z��;���]�a"Rp��'�j���tv����51�$�-�M�<��h8g������]4���4�mU�OC���@��Jh�$�x��0V[����o=�n2ر����Z�n&�,4��f�^�͓F�2��N�{�e=D��-{W^U����~T�������llD: ��IY�������C�x�q�40Nm��Orj8-<a.Ǜ �Xi��[D�\��$c�q��_��ωS���b��c@VH�DpbH�2�(2D,j�(P V �9�=~�{���/{�3:tP��/_�2p\,{�/19�"�Lх��g�.���k�_���c�C�LUD !@�	��"j&�2,{�TV�=�AJ�z^��/V�f�[�z#�aZ��A�W�6�;��|Ǖ읬���x�T���|0�=OY驐��J�>����&r*���ȌUD'����� ���  ��/M"�!H@ \ AB"a��&�a���@գv}S�ɱO}�WVm.��%qk�f�E�x�����
�"X�v	�t��pV��՞���s �7�y��VQ7fQ�GFvkbݧu;&�=��Z2��D�,r�km�6�knH�s�̙��ٶzCR]�i��"��df0��sa��\Z�iֹ�g��֜�,[���.�e��V���	��g��v�99���8n�G bpJ$V�;�\�/b���[����Qa$ ��l�W� �C��"A����fڸ�uU]WWU7�����D�9���%3uWR��U�fD/9����h�!&�#�m��c]����m����˰�g�C�8��4���_�FB�����x--�c氉�e��12W�N�&�-4ZH.���,-�1��0�hp�o<[��N?w���� �痼в��2Ii�^&"!V��`@��bu_<�-�����@r#�V�:����֧Rd��j�Q-�X�ͬ��#F�=k�gL
M���;�͜,����0�~��LI��cM� ��.����U�ί�&W��u�Ĺ����0Ź��:`���RU�����,�F�h�N&5�@���ҋ,��� �Ō��v��-�Ӷ�/��S���9S�˹V��n ���x���q@x��H	���	��Rm"�{I���$7&؎-GZ�-z	��@S7݉�/?\��w�(A�e�><�F����0�-dK�tT����Ͱ�fJ��m=��px�TQo9'i��Oh9��z�H@��9h6��t	�x��"[Ğ�R�[��ڹ^U�:���(DD?�b"!&a�&!������K�4�@�NSUj������F��	3+丮[�^Y�A�6���u��4��%_i<�:>AE#�ŝq�cn�l���l��i���Y6o%�m��z���������ӌl��<���	$ig'�4=�%�y)�T@��;�ʾ�i���!�Q� a3-$�!:�O ��x���$��.�����{�����W{8��Y�#C��ť�q2U����u��[��KXʁ$ih�7rǳ<@������3̃�T
�q	�SS�J�9r&"f�5��������Ƿ���#H�4��{S�e�I �Y�`�u�lXk ��S�p��-&7����d�Ɓ$v��xA��K%f�J�q%�Y6�;�����͇�M�����@�8�@:�}f%���Z[�*z\�<CA�/ނ˰ �d"1�6 a�z�	� >�F���N�!����]���s�x�33SZ��35M�oZXAh1d�v��tD�4wA0Uk�a��j��A���O fS>��������_w>����{�6}t R�(&Ue��r��:�v]�_�oۛ�~w�~ْ���4�F��=����zgK����]R�Rsu�f��S�T_䌒�I�5�9FK��֤����y��۳��K��e1��C;mC����?_���)+��;�-dA��]fu�P�k"E��ܲ��j��=�����4��`��M��C� y��� ��D#8I�(O�I����a+i�K� �a����e==�]a�`�@�����뉭B�3��^5�9=D��u�@�� q��H��!i����ffLI��nf��t�k���wǾ�b��=ɼ)94�2���qҀ.S N�j]{
�DMH���!<�R/�]��<��F�(��G���w�d��d=��O�.Kݛ��w&��/�d=ė�pZ;^k��iԮ�a
&ˇ&�;�ǭH.(kͿ�B�`�7�^��皅�>q�P��5�E�#���p&�'��\e��X��4�7�8c(NU���G�9�z�(+��t|�L§�g��4PNX�M�(n�8���TUQE,�U!HPDR �PP%%DD R-�aD �Hq���<�w=��	%�[ 2~0�U�i���'Jm"�����y᳛6�e�Jh�"����̱$n2���cٞ8�:lŅD�s�K"1�7Ý�#���	�55�9�a9�Y�ݬ':Lb[F\<��	�06g6u�8$̈)˺�.�^'�(����6Xp�]fF�
ض�h`���-ƍ��WcxM�A���`�_��Y
%����l3����`$1b�(�q9�˸��/�%O���M���~޲y��j���uw������8�'U���Lgs	��S��8�ϸ�E��=ztD���d�qrc
I�`�����0H�8��[�+b�n��wA@�e:e-�, ��l�Ĉ]��68"E��ѽ��$#�,�XH��@S3B.��L�\QP�j�s�����+��[��q'� ��zN�VS�c"!�iM����k�,@�<d�u[�
:Y��}y�e��IZ}����w�KbjmMl���1M6�ߏ�m���j�yK6c�:�L�h���ƋO���LJ��F�T�����1��j�k���~��n�|���A�����;I,Œkq�)��:�`x	���=̚�0Zt�U�:\ܦY��� ��C��w��8�T���:����zNpmt��8���_u|߽�.ZR����F1w��6���@H���B��d����!�S��K\�Z[����g��=����� ��wd�9��ÓY�~0Z�P"+}�}�2V^]f�:���Y9}�\���?[�ʃ�UuWW=1�}�v[������ޔ;lV��pc�����+�Uy�-�pJ]�-�˵��K-�1��n���̒����'�-#����aL���Ѧo�F�*֛ O�1�f�4����xK�r���ۓ�o�{O����K�k/!l���<
��� �oe�-���n��;0z���&���n1�|Um9Yͷ2�!���o��liPF��,�F���{u�S'�ܗ_o�OU,P����C�w1� ���y�"n���L�o��� Qhh�\��	�a1C�i�5r:���{(��\=�Ӊk��C����<-��f}��	(f�b�&��p��/u��<��?CƏp@Y&Z6߄�~eLtD�M�M�<�e��� �R�@�:��!E�����|�̋y�f�6�h�I��#�d6�DK���33"I"���xwq
z�3/"[� u��7��ｐ'�^A8�2����q-�Q�
b���O�I=+KI�&Ho�x�+$ c����w�U��X�i*4R*���9�pՄ�d���9�!�s��dD	��P�k�9�s��∂ � ���s�����_�ų��<�._�Dj
���3��ׁ�Q��%�<D]/z�քԺ�FBLaqD�z�$�bL�q	���'�bk�ѻ�9�>�z�SJ�=Va�2*�z�`�x�u颭c��<�N�x������M�r-�� z=wJ�n�-Pzx|�|�ȃ������Da����uV�Bqc�	s/EK&��Ҳ"""!"R��P���f[*aJj�B�EM]�AiKĹ#J�K��FP@j��DLF8v��������/��Ske���`�i5����f��m���`����:,4���5��1�۳by�Չ{Wk�p�HZש����%��,�HJA0�I��j���v&�u�A���[\sv�f2�%�l�����d��6W�[��M�1^:���6���0`�Q㶠�n�n�v̚�N۳WC';yi�������ő��N���m�����<�rq#uR�1�Dv�u�S�7���c���Op��É���a���C@QC<HB��HДRPb4.!�"He��?X��~����\�vݩ	f��F�J�ZVFm��Ubs*����[�2� �sv�����ܻ��ݱ�V��'>�8n���=����)�kp^�0�(ڞI�"�'����e��4�f����i	��m� �\zØ���Qf�}�g�� �����Y���� �M�n��~{>�y7w�NC73V�	m���N9o�
�B��*:�� D77I<R!��"�G�C�P��x0���"�3^���Ǎ�ɶ����7����y7�㖇	Q[��F����[����L��-���e�kl$�u�%�Y��!O*�O(���T���P��V�lm1�+ =���0rt�5� 6��\�{�>s�O��߼��]1,��r͡�"!��	��im6gL���P�m|[�&�}�đn6t?|_��N��F�68�F�4�tݷ���f��w��N{W�2��_?+�̘�^M��s��v�z�jyߩ�|��ʺ~~Á:�	c�'����˖h�KY	���}�Y�ڔ�L�rނA��e�` ������^��W�Ҙ`@A"pH� uz1gNe����$�� H!0��4Sir��V�7F�MD��Z�1n�iY���lҽ`,Q*C�B�H&fr���U4K(�,�6�e�JY�wwq�y���>,%�7�d	��H�{ 9`�og�Kq�:>p<��ؾ!D����츖����Zئ ws�1S2��x��D'��
$i`�p+ N�J��xX1N��QO�EN"Ë�v ��Á>-T����}���i-��.�,-!��+M�8px�"�D<'��Smn�[f|b�f�~�;��[������Ks ���p��fx�T�$��u���{����L�� 0�4�~M ��,�f���g�y Hv�L�����o�m����sy���m���k���|珝�@;�j:r�R���0|h���o�;]#M ŭ�ͬE^������z��i���ԡ6�x� �e�|��uR{Wʼ��E�!�5�����5�x�����[�Q�̘Y�����[Hdu�1�f��6��>.X4��uW<���F�b,��[��<[i-��>�0 " [�f��d^]�~+�ɞwy�}��=�m����o��X ����V�Y�콢n�sp��]�k,��6nE�����BB׺͜HkW`�g�6��l�|���v�ix���/�럞N$0���Ӡ ���d=�<�%���4���w�٦ۘ (<a��� �"囎Z��B���p)`&dB)$���%DDAU"&&��H �����p'� ��0Cѕ�6P��IJ��p� �)s ,��)�-�x
�y���@�+�� �L�D<'�wx�xx):P��'��6�/��;�K<�1kc�6���X9����yͿ���i��T({<�e[�{�]KT�yT��N{Z�U>À��]�S����0���ț�|`gՕ �I�9�Oj�r�L��}�fֻʝ��V��yEo�22|�ˣ�`�맸���VF�D�d�j1F)�����������Ҷ���vgƱ%B(S�)F����t:�q��$�bERMQDPM4�5TUE-)M%DS$E+BD4�+ R�UDąSRQT-,��54�Ĕ��#���<B�@�)0S�=!��U8\�C��p'Ź�6[�s�a��>0�D�H���������L|8�]��$nRt�p�^g�{q<`��!E�p%��T[KS�@���,�q��P�U�r3��>!�Y�oN�UMTJ""Q	8p������e�X�c���4F�@�Vk S�[��|Ƙ�I��p�˲�'�ړh�~w�������N�" �݀��ccm'�S���O��'�N����������	B"�RV�苎K�q^W�7c������Q�!#�2��Ԫ�
���-̘Ŕ�Gm�٘�eѦ�Γl|����������r'�0,�X�d�u�D��*�x�쨑c�ih.ƀ sOO '��i=�ϝv7�-�ClMY[�[+]����${�[7��}�!����=@{R��.�Dd�r�v���|:N��0�� -�\�&���Gt�*�İ〶����[E���R0���C���H� û�a\�
 ����^�{�-F��3�Z���� ��:s�x���U>��~|�Z�o	��D7�#ܫ��ee��� �@H�-��A��֣5�w����}�z�"~�o~�n�@1�4'[�	��XM�6�� x�>b�,w=���ƈS2�I[c�W��P_U��s��;̻C��K..��Iw#_~>�}�?���t�$i�	�E�� ��C���`��2x� ���U�'��&;}_����p6%��@f]��S0�Ӧ&�f�/P-$7�D<DD*( � -W��KYw���i�d��yk�%��b;FE�2iaH,E�]�H�sumW]�������JP��khH�z8��=�n&�"�V�t\/m���Lm�0\��2�a��j,�EQF����c�(2�Ѥ����Yy���5y�4�mo%p���|k�P'���bM�> zA��|�8�w��"(1M���r�GW�\"�WW
���#���Z�\K[$H���]�h�x 'y�������KJ�.����l�{�I�O�	� ��H�vߞkS)W\Ky�;r��t�Ϳ�G��t�<�.���SM%��~��Q]A�����h��.T�}�Ȯ���r&e��f��i�#���p*����1�#�(
��Han���XUs2E��2�VW��w�f��T���"I1%��Yu�s�yqNF�<��<ɗ����&���/�y�q��3Q3[�4��T<�6@�`���.�UD1`e�����-�z����vz�J�y��02^�p*��Ci�Z6�CD<�a[���K�DX� j�!cZ���@��i�Dլh�� DE�&RɉpK�4�B""" C���p��\��� @y���jϱ��-�\���y�e��R�*�[Ǘ���yK����^�p�AF^�(��'=�/q�б�n.����\HŞS�k�y?�9�iz|�&�:U7V�${��}q/rc)T��� �d�P��y�KDe���)��,xR��c��NJ���٫�F�z��^��+1F�TIb�U��wU}�Re�ō�KZ� U-P����i)"��˴�b�H�`�V- �.D�6���'Iήo7"m�W��ǵ�r���v�敧Ul��3Ё7m>$�F庉�=z$���[�oR���7m�8+ ᧑p�ɼ��f�rq�n�t�8@�ݮ^#y݈ݹz��G2�Ӕ�vzMn���)b��.��yX��z4\We-Ñ8� ��x}+a"d�ٸ�6�i�mEuC^Z<�۷]{1/�lV��s#F�/N�N-������d�Mt'�~��G�#��(���;ď|~"��~����M��*ne��䶁�L B"H�&���F���t�[p�,����]=�ƩeJ�"��dsP�荳s��7��
�FdK�ĉJ):�O�:Ї�b3��I�O�Sm� �x#��
���Lu���v�-������2���R��LW��#����;�|�U�mjG�F�@��Rt@7�}��@I�v`p\}���|�ZHDrv��p%��B��>mb`���s�V-2)D����ZZ����pZ`�UQ� D;��OR�WŨ�ce���:��l�5��O����,�z.#PXf�c�ET=�n�g, gUB� �-�p�:���
Z@��tAD�P����$�Pa'�<Xe�Lc��눉oGŬ���o�)�������\��a�e�Vt�Ф���6/c�Y�a���mS���8�bv�4Z"!��4���9��90��kǟ�d>|�|#y��c!'H� ou���(�_8�,rKm�I����uY�������H" �ƒ��ӂYȻP:{$�h�=��%Y�@��ճuz��e�Lp� q<��F�3�B:,)��[֐���ں�I%�8��#��Y�mĚ/ ��(���a����ݶ��j`�dނ&���e�ّں�����xv��#N�ݜ�vw�)D<wm�Yu�Y&��6���}9�<�h&W�Οn;V@�k�4*�Yu�(����fpdss��E��c����ZΖ��Zt��W<�rK�W��_9\�e��Lշff�K�ե������m�<��-�Le�ۼ�@s4��@;�A[V搴��hi�\���˩7������1�Sia����΢���'y�sU���cIy��5�;��m�3kK!����<��t�b�Z���ʀ!����O�a�(L�����*T�3��0~��!��q���ϟ�c�o�]e���:�n������:m�Ш��Z���1��a��d��`��6�[z�%��> Q��Oל��������L�M��閭��L�߮^��%�y��o}y�t���}L0X�W�����:�M�r�9��7e�kG[��Z�\��HJ*���G��튄�z�&��m��c�k��p���<(H���\��Gr�y�5!��gm��i��h6���a.Ǜb�d� ֒awC�<�Ħ�}ݕk:_}�]-��Jݵl�o[v��~���0���[��cG$'�漵��]�]O/\|Ch:���sĺ�E�o695�-�秙����!e�������Oo��~���
�n�b^l��Z�D"!�/�����{-��H�x=��v������X ͧ������O�d���B���dY��O�o�ME獪�&�z�$§{�Q�V�}T���^�Ŝ�z̙�3Sv��O�/�*J�U�/2r��虩uQ��/b��)�/Me�$��YPeVM]�c��o��+TZ��|2��w&�3��+��1L��r�.��J<=���_����ڹ�8Ñ��=��y�T������*-p��tF�o<����]�G�Oq-�Q�1��hB+�5S5f��]0�&+��]>���������>�3� [m��i��F�-0����hMN���u��m��bJ���+�Sj�m{��	��X��� ��$n���Y�����������V����m Y�m$�<@��YI�?T����:CE��5_)�p����>�~/Ѕ�߾��w6�_��yy����g�y؁ꪊ�t��A�"���F�.��Κ�뺖=S		�N;lp v�WR�zE������!���O����b�r��j��,<eә-�5O<�`[�̨��1���BΜ�@Y�$�q�'f��;�t"���"EAp���	;�0�,�"���5�츐7��8�	mo�ԫ˕=R5�31 x�c���n�4�s6`Z�󥤍4ņ�c�m�{u�W[^�w�~�.Z��Iv��Nb �w1��Ì!�ovӰ�\���L��[ŧ�i'��Y9-�tI�D	�``x�.��6�cGKQ�آ1��2%Aw1�B�E:Q^"��jc�,X@�y.�:|<-��r�y�C, d�����6t�o8���L=��06�34�����1a�=��
2&D��ƌ��3W���<���{uۀi�g��5t��YϛU�$i⧔�� \qlv�}�t�	CM��Q�� �D���ɗ}^L�+6~f�����7����E���k�z�u!�����t+9ђx�k�:�pk�cwlm�"Đ�	��b�M�L�~8�|�v��sRsE�hf��9opT��f�86'K�w"
�q<`�����&�8݅���o�OuÉ�-6e�r�P $�B��!�<�!)4�L̳sc�(#�A�!O�p"BYpޘ��x�4� ��g�| 2ǈ��mq�,$��a�Aޥ#��-�-�uЎfXH�D$��AE���ܹQM���������Q�e�X���\HEuH#��gi�N�z�E�e\�����M=-����x�8�؞�O��3Q�a�T��Bu,�iI.�c����C�����B�;v�#�M������Ì0���y�������mc���A�ڋx�-�d=�Ӊ<t��掵vC�U,K]������VN�mrq����� 6�%߲a����0h�~S�@�6ܚ�h��69Ya�4�~�e��w9Y���_l�>�Cn0�H��R�$K-/n� �����@��X�"XЁ1���)���5d
Z1,��J��C�:E�#Q	�1�Baӌ!X�m�EB񘈉���C�zS8����c��C�D��3tC�a���S��9�h��ޕ/S�w���ڀ�<=3b̌8.5��d>TO��Ǯ^Ӫ��!�����<�5�x@�T�YT��y�3��M�Sr�9wR���Yy�W�=�F�	����ǉǙC*#3諌��I%�s����5`EH���m�E@B� "ha�jX���#�K�j �^��[a��] �3����穄\�E;bڇ\�`���u��xBn;�x��m���5!F�=�p�g��v�A����k�������R���5�lW܊f"�릊�8�6�u��^q��6ܲK}����$b�F�U� ���\���۷7���x�dǩ�e�bx�e�l�B�6Q`���hp�v�s���y �d�j�F]:��z{�QGN�:mI3���`��(( ��|�Q����+�"�"�=�_�����7\�m��6@����9/��*T�W�U���s;$N��.�����`}�ɵ���]�=q�����o¾w'z��뺯z��@=v�Js]���`�<?�Y�i��Ґ4�c� [b��\�H`��Gs�D��|k�@O��������p��W sA�T����y��Y�%�׷�%Nꯪ:۷�Ӥ�D$�$sf!�&�}��G��9�o� EÍx�����s:a�o�{q<nSx�>��D	;L�ڲ�6���8m�=����^�Z���*����)��a��!{c�0��z�,���s�eC���b����(��y�~p,�����N�ƦL5�߯��}��y��S6鬷Ke�.f��x4 ��R[�o=ˑ�1o1�!1�Z�T��1��a��zyNa�^ �O#�{3�B_�X��~�F�װn�nְo���~-�vD�UUP�ܗxN]D	BP!�"�K#���ό@��� 'qA QF4�[�Ζ|�l[�	�}m�4�4ů4od<���a����,h�C1]�˻�����w�'~�#;Oپ��W|�
F�� �.�����ήH	c:!u��v�n�ֱ������ZW��I��u��`�y�n.�z��+���v�PgsRv�0Zȓ�	���`��Ȳg K��&V�8��`^.GV�RáQ���onr��Xgv��01��bDn���ͅ�˒��_u���+�y�K{PA#2��Q鞟ey��E����x��E�q�N�����m�y�h4��~�����ޟ/��3x�n^���1 ���� ��z��]�!�-4�U�WP◖��xɧ7=C��u��4=P�knI�[ h�W�7+���?f��	|�æ���-ql���&1�/�}���+��]�^�f�z��U�Uû��n��lo⏮��`�\x٧��^��������<#$�>v4Z]���Y1��u����祉��K�c
h�+dB�YZ)��7����m��f����ioB�ʓ������
A&F�~�Y��｝~����oY��u����o��RZ�US�����������\PE�4c����{��<����X ;x����:��,7SE�l������ƙ]�S��1�WT^��6@bCH�UץX���i<m��XE��8��u_>�5m�f�W��__�τu�N���Y�M��c)w9��>����G��f�i�O��Y�8���mh[ώ.�r���n�;����� !����26T��O.�:+�"��7����g���c��a�-ʱlH��W��R%���fz�g����A#hR�~�����i���O�ފ7e]*h|V-Z�g���C,�G�su{�ڈ�7���&Ǟi�"�>���)��'���5oM���5�(E������p�r���	19j+)�<�+�{���J>QUk�yUG�"�_f��Tn��Uh�T�T�ɧJrI;�B�&X�Ia;��H?�(�/
���g���F; T�"�T8�C�$�(h)+�DD�Q0DRL3LLĒM0A$�1KMC2�0�A�Ib0�#$�L�K�I&0ቂX�d��B	�$0LD�$$D���0���!��c�QBLPL�%2"C�&3��y�ƾQ����K]@�<��v	�uCt ����,�,�C3+s�u_��\�T�S��{ ����s�E�[y�[-bz��5F���]:�'K��e�rsbQ���>�M z;�{@`Po�_|F0I�ʇV2��]�˵ĝ-�>}����O>R�y�/SC��\��|�`x-��Ctߡ�Z���S�lv:�� (fm�����L���{��ݾ��߽�s�n�λ���WS�t���i�y�����l@�&�q�0�Uz�3cg�۶�ϼ+�27��u^�]q�]t�]`G��~~����h$��z冶0�Z'Vr�� *#G��ه5c@��g�y+�b�	��or|�*�������[v��^쵍l��i�ǝ��|�/$�QXv'Y*�>=��W�	�� � ��,�`�`s�E�����ï�/N3o��'��ud���Y��b^h�iai<DCòw��Vـ��Է�s iCm�!�
��!%( oݚבx+�n;��ȯxz�U�[Ň�lð� M���}]�����t����|��*]��6��) ���rw�����\�[���P����6����50�:� ø��1q������wc�E: ʧ�x�Ӓ=�l*faDND@�pC�B�ey��� �G?�j�vE��w�t5�X�\�{�����Q��:�]W��_HK��1	�d]l"���ܜC.d�)QBf|�We�\�_97�RA
D	�h��p���z�S��i݉���#;�	lR�Bi NM)��M1�0�q�%�ɀe��x�A9�K�DL�$�̩��.N�<�l��(`����/�އa�l:�-U����ɽ�����Z�uG� ��*1�֦MF^^]����ܓ����zktQH��W"��xt"M�6w��ꗎ͆徸��Dn���X�9���zx�]p�`	�d�p�p T�xc]-�A�s$��������h�*��W��kx�á����0�/�"���ۯE��x��1oό�\��u�ګaͬ,��1O2�wx)ч0�A*A"=>��)N�s���֦vZO~v�ެ����b�,PD �Θ�f؉�Z�;ٻ���M朋p/��}~ێ�l32�br�]C�xx��J!�m���d�]��sXh�f���n7�A���x-L0���C��tφ�׆ޠ�<��q�pd`��g�z�������UUSUUUUR�d�  �D�_�>�P~.=����e+��#,�R{�ә3������&�v�!s�Pf�&��}A�׻0�N��4��:��!&�I!Μ		����ML�7	p�zݐ!��@�M�	a FC� �`p�VH	(����� �"D2���
`�(W�
�u8	޽+��RprD��0H��P�@ e8�U5��\��
���AXEt��-�P��E�,*� !�� g �r��"e &R"i� #�"$"�@P�H�Fq(!��{�w"�!a�S��^���0����`,�p6�N0�]�\ć�8Hb��@�檪���ENo��H�R�EB�)UE(��*!y��y�9Vx�̛�N���.|M�sq���<�p98�a:�?�6ן#���%~_��g&�6�$�����Fw���v:�$ř��9�Pu��\��״G����f��@O\!��Oo9Å�~�԰DUO)��~}?�g�a}�8�����,>����=�s|��H�>=X���w�K��������{� ��@I""�~c��I�(
� {�?���:u���x]_R�N�������?��e� h�o�A�Q���N�^Ԍ��s(Fi��9�x�=G�p4 �U5�"�#R�����=oü}�&��c���|	�(>�s֚;��	��ҟ!!�~��!|>/!!tCÒ_���2� kX��A�G���� �?�,;��BrN��3���~��9�?��#�0� 򫋇ߐo�����x#�9�<s6� ̌�0�^�r�S���L, �U�c�����=���L3$޽��I�E$� �C�`��!
��6Vr��@bV D�caA
��*
�T1	@ЍHP�I�� C���#,��H!@B,2 �0(RJҴ% �0ʂ���ʈ2�K*0��
�"K-K�21,�&�08e&ZV 
&h�3$UP��H �$ LH��Mߠ`�	&��@/���O�>�C�@!N�2Oq�1�oxO�.ܙ����O����v��oSp(:�w�(P Yf��n:}�t�=>9�'j� �n�L2�	�t�6� �\BX,��=+�9�w��)	��D�8�����#��	�z�;�r��P�G�S��4�����}�rk�x}_���ة����a��s7�a��	\>RP�QCICICIICIHRRP�P��P�RL�RP�R�RR�D��RP�P�P��RQIICCC@P��P�K,KKICIIE%CI0Ĕ%$��P��0�K,4%%��4�1%%%%)IICKCIICIIM��3%%%%%IICICIJL�����CIKII CIIE%�L4�%%$DI	$CICIICICE%,��AIICI$�RRP�%$�C2D�RD1$KIICIIE%%�C4�4����4�1%CQE$��$CI2P�RPRRL-%%-IIE%-%-%%%-�%%%-%%!ICCICBP�IICICICCII1IICI@P��4��RRPĴ�ICIIM%$@RP�RD4��RR�#I�%%	II12D�4�4�44�%2HP�P�RP�%DKCIKCICIILIKKICIICKIRR�P�IC44L��4���4�44C%%-%%E%%-KICKIE%$CC�R���1%IICIKQCPĔIICIIA2D�4�4�4��%��%-%%$CDIICIC2Д1%%%%CKI�Ĕ4RҔ1%%%%%%$CI�RR�RQ0Ҕ�R�KCCIE$�CI��1IIM%-%%D�%%$C���P�IICCCIC��4RL��@RP��RRP�P���44%$E%%%%-��4�-%%-$IE-$CICICC0�QRPĴ�%%II�D4�4��%��441-%ICE�CC�RP�ĔRP���4�4��4R�44����1%$E$ICI�Ĕ4��P�L��4��4�-�%$CIKCICE$ICICCC�ĔP�R1$KIC�P�II41)ICICD,�CCC0�P�CI�R��P�D���44�4�CCCAIICP�T4�D�EQEEE1QMSTD�E$EQALQAMB�-%$y���� ���b�I�l�)��#��;��`?��tO�b	֘�ya7����_�#������>��)�#c���#4�:�r�P~���Y/V<���&�RO{���ǥ;\�#��6ӷ�&���%/�=���1��=����<��Ǵw}$���悪�Ν�k	�M��9�Ф}c�@���6���s��k��`A���9f8YrR${��<�o�f!���M����,��nE@F�j}�y�}��C�aC��4�����Z4�L	���o��L'�oL���S�Y� tՄ5x�.���A��M1�Jj442`�Oa�}�ֺ�`4Xs�rN�
�
���!3EH����l>>�66��@8�2O�pt'$�9��2`8�H�!���?�z��oEw��e9i�30�8�,��߿x��@�a<Na���{�zO^8L�$p3� ��sa&0	��*�	2�c�����q��q���0(������� ��w�p� H��!�My��#�"?���q�����}3������u���N� 1��0^��5;�B��&���	���r}G�����6)�I�Ϙ�!��G��y$9az?:@�<�C�f`�
�ztO�ޟ�ws�v��'x�U��i=HzOq�^
(�L�b��00�)���D`=h���T�O�EMA:d�o���S����7�^�P:MX�y����ϲ�h��8᪚�+ CI"A���̳�ޅ���D�1F��|�L'�	b/p~�>�����$�7'�@���y�y��<�M��(E�9���pJn �錃�7o�y�̰�l��⪮�K�:4��|w�MƦ�*���;��"3����x���|%!R����^<����6_̆�3� }P�2i׼D����7<��{3�;��s'�����!9�
j��a}c�C08�8�؛�	ڛ�9�Q\�b'�r���1���s�9�ࢀ�Q��?_�0<;�"�UA��a0�}bh'�3�� � � I2#��ܻ�����C� �;��x	�6��xfz��: eȍ���;��/�4���0?�ǀ�=�:�yVA�7hg����9�_��f�A/��!�c@6��U��rE8P��([8