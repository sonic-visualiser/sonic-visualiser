BZh91AY&SY�@���߀ryg����������`��}	       p@        �|��EB��B�UET+ =�%��6���������k��LܹGM�˔(��yb� gX�E�(Cvu��5w\Q@)պ� �Q��ܠSW;�(�8 !�@�㛗�QG7.(�B�nX��x>��s@(\�(�4)� ��Os:�GG@gr�
(�W;���GM[�QE:��Q�EÔ�듼Q�@�t�QA��  /GMo,@U[�(��易N� ��          :�   4�	���@��ha �  �LTT�� 4  �L�  O2���*dM 44�40�Ȩ�%OS  L�` & C	���I*h4i�@      E&�	�i�4i��*l�����OH�M�(�)��OO�z����nt�$A|�C�J&�6�"D�BHC�7"%?��sp	Вj?�������^�n_������ڕ�a�_�-����~Y�O�8����wX����I�U�x�I���{;�D���tTsڽ�KF��ն�ѿ����R�I$*�z p�)]*y�wk]U��=\ڋ���u���[�{>eշd��D�B~��M؞V���g���G�5ӿ�������G��wU���������������|�M��fo{��3FS,e2ť��iY������\�Rش�z2�dQ]N(�E(������~qEq���ݮ�+�R�تe��͙�2�S,[s8336e��͙�����e�KN.S8�ٖ2�ť���c)im��2�RԪffl����Z[�ť��iis37��y���.gX�e-��S{ռ3F��c)le--�KL����ilj�33{�3Q��[iilZZ��L�ii��ffl���ff̦X�e8���X�[�����]S�kL����2���S)m������3322��c)��꘦X�-KKh�EwqE(Ӝ���ҙN.R���qc)�2�R�.^)���X�e��S,e2�kYL�ffo{�FS,e33�38��SW)����ʙL�X�fg[���S,e2�f���FRӎ8�)sFff�)lfh�e�ffa�5uL�X���L���qr�Kbӆj333xe-��R�KKb�ʙL�X�e.j�ҳQ��---�J�\�q�������2�c)����L���--��X��e����4fffc)�2��ťfpj�f�{����{���ᙜb�*b�L���\ե�{l�ʜ�r�*e�f��]STŌ�fqKKc��MS,e35K�2�R���e8���,b�R��e�\�S,V�e��)lfj2���f��le���c3FSZ���{�n���n�c)��Lf��]X��M�qKKc)���8���ilZU8�Q���)��L�ii�2��)��8���љ���,e2��e-��X�fh��cWY�����2�b����e.g��lZe�L�X�~4��h�噽�L��������FX�є��2�c)�1L�b�)sV����--��)�2���kT�Ռ�X��b�,j�2�cje��X�L��KL��ڦS3FX��\��
qN,fh��S3S�W*r���NV7L���e��bܦS,e1c)�Ō�S-f�����L�b���i�����i��L�S-S)�2�c)��4e2�e2�)�1c)�2�cw/ӌ���X�e2�,e2�b�S3FX�[���Sw5�bشʙ���X��n�5L����S,e2�\�R�e2�S)�2�����e��,e+4e��)nS)�2�c�2�)���֎T�˖f����T��і2���L�f���������-����xfhŌ�X�e2�S,n�s�Mش��c4e2ŦS�8���b�,c5Kc3FX���锶--���n�wX�F�qE;��߷`  �S���ʜ\���2��Y��~W�0�I�~��ƪ��a?���W���&!Ῠ���'�'�?�A��~�!��7�6��>�݅�H`�H!i�ȵ����S��L�Ur���b��/RqŽ;�\�[��!�Z�������q�p:��(�ND�QhX�i�bLC�A�y\��6.TA�xi�q�8�a��a���Lࡈ%# �Ub�!H���s�6mN5<(�pq旦��'�N��;��,�ߓ������T�D��3Ys�|>%J������&��ZBp�c�<I�\T�]��x���\:2�
�F̉�G���H�����X{��O�)S����#$Ma��� ��r��Y��AO:���rni��%�T�9R�U3%cҕT��Rǹ"o$Ҁ�	��D��ˉ�K۵�xe�/v�*���$�xC����5534}O�82�)����*.p�u7������d�FC̡����ɉ�z"�2�*�70,Qi���٨�&#�Yu#���a�U���E�M�ý���M=�P\�M)S�T08|S9$����⻔J��^���R�r`�`͕St�"%�\E��&-F��)�
���d�T)zy���Z��i�ʋ�N�ndN<'�w�� ɛ��)K�Z͹0he�{8(S�����̘��-X�n�E�Jrd�*���Lq�>`��v����+�-N�S���jhA������6�@7V��8BE�
C�
����V9�/u*��{��B��lo9�O��SAZ7s�8�Ÿ/�)���7�$���"��F�䫻�o���,Ud��ܹP�.�'#,Q�Y"�]5Q��/��b����j�TB�	�@�"`�Qj30UE:�R*��#� �v���!�(TJI�Ⱜ��ȩ���fe>W�ȉ5$r2�t��UV-�r����1B�5K-eLL�sb�Y|���5X˚z��p�6�ȁiR��S�fC�A�B�8yi�1�P/Sxd��as/��UX.�2�I8`Ҋky�w6��1���
�"�<�!pU,�ӶTԊ�I����a�I�Ǽ���zz�y��9�ˈ��zJ	4I����yy*# \�uc*���$�x�����-�?��f)������[�y0a9D�2.�UYk�{��J��8c��iB�(ׅ�M�\^E�˪����-�ẇPR��B"�M��+�+E]�9v��Yz��R�̗�x9��S�R��Mڻ��ܧ��q�A�e��*���Ud*�{�J��zx��5�B�2�����2)@��2TPɜ�|&K��M���Y��Dc�PBk%��wFP�f%�r�]۹��B�6�]������𨜘�ʪs�B�ڷ�������nl@�����r�T��E������'*M<�ʅ+&*1�Xx0�z�מl)�E)�r�5s�Ys.�Ș�Ǣ�)��5�IC/*a�2&�#j��9��B��EE�B�
H�4�����*�\��E�).s2�r'3"S<ନ�0�`�]�̼�Y0(��N.DCع2*��a�B�T�A��7���!!99Ys@�vM�LK��.�/v��Rf�#D�e�O��7J��Ĝ�x�6חT��H�Yd����g�V��ӂ�<b( �n��X*�<U,|�u&���TL]�yǃ3Oq	��c�U_����?`�����߮J�ܩ���R�!U�U # @�q�tI�-M	0�PK�H  �`)[�� ��4 H��
B�� Pݩ��  j�Q �-
P�+*b@�ՐU Av��IH  
%m��� ��C%n䩷"�X� ���Z! @"��� �]� 2ɠX��,h@"�P.�d RHƂ۔����(�p5pP3
�@@L��M8��
n� ��6,M X�e�$ ���.�E�f��4�  � �@�!Wu"�\@���� ������>��W�un���>�W��3m�/�~��ӷ�۪�;�g_g��ǫ�Ý�8��^<<��˽�:[���N|K#V�3���
��;���#��Y?R�ѽ�]��g�7�W�瞿4?W���5��0*:���)rQK�n�5u��f�r����L[v ۍ�D F�o��R.SL:	��e��Ɍ�A��ب������)"C����].m!�^�aէw۟)���Bm:�i�Vء�+4eR�<�\��s��Jp��A6�R�1����m���R*�,��al ][�$z�lJA�m���f.xQ���TՂ�nJf�9�
��X�*�X䃳�7jBc�ff��d�Ѷ��l�F���d&r	a�̘3Wl%���T�lM�wv��a��8�9�]���5��Z�֦�n���:%a���II�tR.`P���nL+i�ЎWWV�ve�&��
,�j�U��˻s�I�D<��[6�M�1-1 ݘ�
MF457ICnjB9���
���n�)߄��<�պ,&�4M��V&
�y�-HY)�4�,���1�g��-rʬ��CP��F�5�Ú�l����[Q�.��������%����른m�Ѥͺ��g�86Q��12Q��hXfm��\��]l4Gf�lQ%"y��{B�x�m���f�\��
R&̪����6J<�-!,c�E�n��ō�Jn)�ݺe-U�k`�%O;ǭl�GA�c��e��fW&6`�"�KpLgh��R0r��e�Xm�V�xh鮘���aL�Csl�M��5`���2����cju+&��D� R�j�`^����5|� ��`�qa����fB3R��k�F�i��1�� �iE���fբL[Ђ����(�mM�EKYc	uճj��7(JD�	e#���2R�U���S��Jl�Δ34W� �]nd��S �; gd��(D�7�u-I[�[�l�Q��E�q�u2�@ M��TU�].%q��Xiu[���U, c��9F&af�����*4�qwk�WT����#�T�,��;��l`�e�$]&!���k4)E�\�l�CdB��a�S��J�����Fպ\�15��掠�\3Z�h	v�6t�+,k�������SnLXM�ؙ��\�ń�b�4y]a5&[.HL����1\xy��q����z7�ם��"HD�Y�=[�]=؞�����"H�<�{���_g���ˬ�H�#�ξ��i�H�fz��<�G�!=�O�}�:������{=H��[��Z���<j]�����b�Ez����ᝎ��A��:K+;��z�<�C�^x$��q�<��l� ���#F�H�+$�<�6�I�Y�=ou^����e���I���Ou/o�C��	�G�~>��u��)m��OH�+	<#g�_,积��������#%bOc��!<m��#<�!�x;==���a�1�G�+!0����\KD8�=�RD��n��8���~%�O�0����Z^n�$���H�VP&�a<�yy~e���>t}���!e��k�C��u���a���{�f�0�be�M���xKd@	���,��Ye��=%�=�Fߟ�>�y�'��Tw���6%&�-)2M�t���f!�d��Zv�ҴgS�l���o��׾[燭�71$�����.g� yt�"ܠ�/$=סZ&-jdVe=<!�fQzx�,P�P���M(!̻���e*��kfB�A�"B*��w񇔜*|��Ͼ��e�ď�?F���s�=��_��4�1����{�ɻ��Q�N$��)�deHp����/$A��R*�|��,�<y2�����{$���)�{����Cn$�60=>����
�'xMg����'|��g��W����<:�z�|���M���,�$ C�˯DT��t�=�u18���:�CǛ<||
}m|�=�T��=3ڧ�=z�C�ӯ
�iRH��O`�������B��9��᷀��%�eW�<��
s"�JH{HѬ)C��PEK��<|Ͼ!}m#(��>}V|��@� F����CD�L�y>����TS�,��.%����go���]zI�kf�s-	��$	3SLn��@�d�����7�+�j�=�Ӌw�M�������@+����ޟ$�	s/�n�]��� PTL&r1C�Zǜ�=��Ԗ�@_oD�'�{�i��>����Εx��cE��W���.��r�n�k8���b*���4֡���u�t� ��5&��9XF���2@�j�3=��U��)��zˬ��O�l���gpI3�;�N�K��ϓ���|8�f�zA�:t����1ӽ;��p�Jwxz3��&`�6�#�1-d
"H
�hxw�)&:S�G2�9�Y��3��e��zq���v��v'�D�
�E�m�>_�7���_&�*;�>��N�o��O�͐�(�f�e�4 ��E��Z]��E�B �0R�7AH�  �L2 �(&�*5`�6�2n��uu\��Ue��g�s��"�)CVT�@T�Bj� b2J�
 !K)��U��6^�A�!YU܉""�7y��\w����Iu�o/���;Elڤk���.4]���\M(#\<��(]�m�!�mi*��D�$Bl9l\�Qc�;@m�9��XVS�qB�;f��Y��@a  YLb؄)F͸��l'J;���U4�d,i�R&lC	��..�5P4�Yn��M�m2�UF#� 63d͵��b*��Z�#fK��Q,�/`pmJ]Pi��Ų��;,���R�-����f]���O~}kv��Z���-�[]5�6�[b֍Qm�smƍƻM�XwU��H��{b�'����◲T�oʬ"�V�٠&f\���lV)��Swv0���E�c�v]�68an[`��a��j�d�,͚4)����(sS9��Y:fmI
��h�R���'�$�;����|�n��2���*����@y��g�i����z>�-�Ky�6m옰��e�aµ ʂ+'8l;���ϓ�z@����n. �т&�����f
H9�Пf�׃v�PF� ���5�����a��lm�L��C����!D<�D!�L���jm�*}v�, �����n5�Ƃ��
^�d�\\E+�!��݅��g`15� +q��T��;�^UuUy�����[oZ�"
A�)Cðֆ��^���ڽn�&�V�45�D�*נ�k�q!F�9�b2��
�Lk��f�ƺ��l�Z9�u��5�-��	�#~?-���!��/XXSh�P��G���X<v�(W���m`6�\0�`��^�� H(E �w�͗n>d�:���1㋙�9�瓮|�'9�*�Rf6�T��pAE�,�m��:[3����B�[<��d�J9�M+l�Vp��c�n��g]v�}>�a@wauö�U��n��Sz����٩���vi�$A[n6�>�3\>��6h��ʹ����2�m2�l��:7mގ�滤�}�2bAȽ�v]�@	�6π�v�����^p� o��y��[�9;�LX^@��!����1��ֵ[�v类�ߞr���Y�|�l/KT� ��	|x�]��-.�h��kDd�k?�v��t��/�������n���:��fY� X:O��l3y��[޶�v������7��zw\
mg�α�(���<,��F2f�H�>*i��3�}�l`S���@k��h��ݕ$�����n�z;m[Noz���zZ�
�A,k^U0���}^a`Kx
��g�b2 DCV$�
A�g���n���]��ۋ����}s��U8�S�wϐ+��ZEV1���:�U0Tl�ݵ���K`�<|���J"0�B!dl��d�"�e��:t�M$[9����&�b�b�	<@}�Ƃ�����,��i�1�ik�ئm�	���oKy������j=c�~z���|l�9�;���	��irdT'������N�}va������0��}T.�e\����ꢢ�U��I`��, 	 0��֚��צL[��v�7ga�ƘKm��'��l�Xs�{��jk��$�-2$� �a� kۍ��vd��ہ� g����⿾���ΓJYѬ�Q�.���G1�fW�I,{
.2�
��@۹)[�H�|��>?��KȺ���Eÿ�O�R\���MM���؂Ϟ���|�;�E+�k�3�����~ ��P�S�N^��b��h�*Mm���}`� ����7�d�Ǫ��R���iU�!�� i�q!���b ���뮺�\���f�m���Fń\��Ԓ��z3����$�#��Y� �7&�q�c1�������/�3�ii#N6[��\<�` 5�C���8�6i���c�ͳ��ض�><�U�� U~�zyÞ�&���"��理��y��n>A�e2&@s�<:x�"	pK�����D,iP��)��VgKa�7w�*���k3+b�v`j�4� 3��V�?�Ky����}���Bƀcny�/�Q�z]n��]N{��"�P� D+�`֯�:2�vK�8�&�؆�ƚ4����)Vb���0S�
A�����s��B��l� �]�`��+��<C�p��@VxG�d8�;�x:Y��0.���x2��V>�A���`��Ţ�[�us�i� e�Ӈ�Q�C�r^��vMh����!����M2wn�6�T<�p�!2��!J�z�8	#i�t�~�:d�8ّ���6 4�l�2.�����dq�v�=Y����$��{
���D%�IO
�Ƙ�-�_���Ȉ�8�NC/=��OwĎ�~���_�a�Ǽ�o[Vũ�3��i' <Z��#�%<��D4�lu����$�;���@1�O�0�=��v�ɨ���揭��q�d����v޾p( ���Qf�&
�q6ܤ���5(;8�FD���4<���Y&�ވil �XD�t�|���`��RB @�P�@NT:��+O���e��߳�D7́����a�d+��i6�,�H��7̨�X�-*�K�!�Zd���5�W>��A� ��N�%�y�w�eQ91V����"DC��s��r�_��;�`�91r8�^d�"�
�07,e��e���'�� �4�^1mU��V,kLk�VZ�.�%<@��-�>lr$8��i}�)n�
��2�7��KYo�q���Q�z��-�t�U�ql��.XmH��9.��b)����	)A9���i��F��ΐ@tIǸ�y����U�h �0��3�n�<	"-���q0U�q��j,6�]��O1ʧH���#���L%�x@hf��	<��gl��I�'Ϟ��y� Z�8c�H�w��Y��=D��r�.Ӱ�)8^sݓ�5J^�����l"?sҟd����l��7\���4����������y�pCԎ�[dkx4Yh	M���
�q`1֭�-�[� <־���B68��e���dѾ���S���OQ-�xZű��s�`Tđ�\������<D�'��H��w �>4}��{�(,����p;o�{�Q�x�i�	v<����L5��$J��a sh�>d��Uw�?=%LJ`Pf��҄E� MX  ED]��#�4�0��� @�!@ MX��\��|o=���Ws	t�w�^�fd�X�� ^bs�E\����φ]��;��ؿy����>�nxs�.%�e��q��!��wr�|u;�ʊ��"G��)Q��K����,�~�y�Dy�+Q��6j��ԇy{�򽓵��0/ꙟ>To�g���=52؉U����C=!�<$�EV��9��������8 R H �B��4P� �!  5p���RX���V���e���*\�uXLVB�����ne��\ �c79KvJ:!,����-"ڣ��a�x��y�]�2�	��rd`����R�-5U��B\ĭsm��ն[V+�)A��%1(���f�[F�&u��-ٖ�u4@eX"��	(0n+���`
V�����cRĶ4�8�+�l�[tX���U�*U,���ZҲ��L1�+\�QK��[ͥ��X1	s��FP�� �>`�,0��~���؈1�D �6-y\ͮ8�EUb�b��亙�Li@ؤb	�%��!��Z���!�	�m\�.������c��^r�x�+6([�\(�d�"��x�1�7�5~��(���ׂ�߆>k��k�Zs%~1��l2�E���� ���`{�	�9v�ŰZd�a�߿��Y$���9�C�ݶ��,B�c,���0+.<��yZ#O����G,��uE�]�O�N��m����e�-l���4m�і�Vt���k��<��Z�6��=L#���S`'���n��ww��9�.s~|�_/��^��#��A�6��7]s��r�\%X������dB7+FZq1��<�(��A|B�Xʾ�a<	"�];i���˓��'r����A�����q@x��H	���	��Rm"�{I���$7&��j:�A����nd1�}ؙ�����p�1�&^C�ϴi�k..Q���D��A��L����l-6������O$>�����󧀴��Rݽp� Kk�Z���<h��-�Ou�n8��X��W�W�q�EJ�!8L|��^�b.~�ʡ/�� ���*������#|�L�9n�F�Z4]�WMl	�Xlg4�X������'V�PmV*�諗	t����Q {�Y��%��cgX�1殞@I#K9>a��, ��O<���� m��&U�;O@7�8D�߱���{�7m�c��e����Im�l]���	�#�
��f��qu"�&B�ť�q2U����u��[��KXʁ$ih�7rǳ<@���b}����<�=#��V�8P������<;��Y �����adi &���ju��z���fW� �ذ�������4Z<LoA���ɵ�H��� ���DBNRx	;�t� �%��ӬY��i���8Z�����1-�U���gX�S������9e�g���n^� �2��>>hC�g����ffD���q��x��|���/����v��tD�4wA0Uk�a��j��A���H��a����ܼ�e�cw=�����M�� �
�� AD�$(;��N����;��Dd��^/q�ո��3�D��F։��O��� <V�`�An؂m��X���h��c��������	 �?q)+��;�-f�r�3�Z�6�Y,��唦�U4����<��[�EM��C�"~sn�� KVd�����-��4V���$��eW�zz+�>�ô�C%�2��e���,��u*���Z�:Š`	��8��$il��}Y:O�>���{�͵�"�2�u]�DC֗tKa�.�{��ܛӐO+�G-(6�j][*�DMH���!<�R/�]��<��F�(��G���w�d��d=��O�.Kݛ��w&��/�d=ė�pZ;^k��iԮ�a
&ˇ&�;�ǭH.(kͿ�B�`�7�^��皅�>q�P��5�E�#���p&�'��\e��X��4�7�8c(NU���G�9�z�(+��t|�L§<�+���Wk^���Z�V�����,j5��,[��(�Jjƨ�ŷ��ַ��1�N����۫m��l ���Ya柹��p��))[��q��{���a�#��Y($�I���I�G�H=�fx�,�I>��DcLZ�s��p~��6��4�7�'>"5!{���I�-�#.m�Pd�_W��w�f�w�����D� �
��t�a�au���m �$�ѷ�[����$���AXņO��,��FZX6��e��DD@�d������e�\���ĩ�׽I��<p��'��� B]��u�U��	԰q��6�a�1�:���f�]mee˘�j	i���0�iV�쬎�g�x_�|�z��띧q���S�R�y���6�a�H���|"�ik��$8!i�<������d�国�::�`sv+@Q�W1�	��ϴ�%w�Kq��$�D!I�
�x�DAi�S��y�� K2t:�\�-܅,�<Ų�h$�->��l��Zb�"D8�t�^�(�
"i�p+2�ګ�@�͆���4�\�48�i��	�$ĬNoUM �����1~�5L���}U�	��7
a�x� fD�
J&��3��W�|���O\���<��G��A�fN�J��K�,4�[�L.�v�n�19G�.a��E����6ޓ�F]>��#e7c/�:0!�QR��mɗ����yK������L�|�{Am"�-�X����ƀ$� <�����0' ��&Y�W�K�{����� �Y� ��>����Y:QW�$ک7���=)X  Blk-6��j�&�.I6��j��ݡb��\�զ  ��t����z.�X�`ԌW���b�xe��4ZGo=��8���L�<� U�6@�cxͱ�A�k!ǁ4���:@���fDȁtQ�E�mќp�>��,�9=�z��oe�-���n��;0z���&���n1�|Um9Y͎elCk��ߝ��Ҡ� τj�y��A6n~�Y�W���!�P�I�9߼�Ķ�+=��F�H�A��v���� �`f8v�CW#�`�����%�޽8���Q Qv���b��[}^�<��]��1`�,�ey�`K3˼�"Əp@Y&Z6߄�lv�:	"�&Ѧ�xѲ�p��{)K K ��(��~�O�Y�o!�m m�� �jG�oDK���33"I"���xwq
z�3/"[� u��o1��{ OƼ� q�e?���[H���i-ԟ��zV���L���p�:p3�"yr|��i������W+\05c1���H�P� ��% � AdD	��P �DA Z� j� �ڗs�3�;�� �PW�n�ê��A��z�E?��	|OKާ��5.�Q�P�\Q1F���<X�S>�\B{x�	����4n��qO�޲�ҸOE՘r������X*�1]zh�X���!S�#=�w�SeÜ�z���]Ҩ���T�"�"2 ⧪>�s�m�*n�U�P�X��\��R𦉨y�����"BD�$
�%��̶Tՠ�P���( �җ�rF�Z�X���ՠ	�������fO�n��.z�H����AeS-�\ˮ�����A����b�L�tt����nBU���v]Wݵ����Q��":�^�1��Е]
m�,fl������0Z�ї@��Kmڸ�)cJˢJ�UB�ۡ��;s6�n,�b�d��Ykce�Lˠ4
���[e�B���r�¡,7\�g��f�0\yJ�+��2a��Z:��T����H��ߟ�	��I���l�ٸ�bMQF�1b�,���m��X�F��Z�X��ލj��Ҷ�!�˗<��~s�_�5 Ւ�R�UK�ҡ��U��nU��-#�scu� �lM����l�Yd�� #�*9�V^c�s-�N��׋[6x�
���U����ӝe��4�f���F��Ƙ�[m�"W�0�0lrY�{!��(-�j3w��K71�@`�4���h��d������E�Eo�rIu�v\N�$����i �߾���$�H��|�y=�B��À6@s`�l�{3��G6&��3�2�x����c���4�`�
:l��h1ΊOЌl�5��;�O�������,��u�%�Y��!O*�O(��LEHLm@��o�mf��b�� �ؽ,�!gKCZ�o�%��������,����mmʊ�I;�|-��锷�t�Jm�/�w��ϡ����#�·��!����Hܗ��gh��.���������{v�|!�g��ߢ�2�E�C�V8���*�q-�IZO��^�p'X�,|d��|�rÍ �k!7��O�k;[R�I�.[�H4���, �3YN�[��
a�E͗s��{�o���>|���y�홿1�! �LD�.<Q^'.�j�Y��j�2���e��	v�5$��6���r0dA�k�`Ǻwؑ��X����O<��=��t�h)�8���� ���,4��<�5�'�� n���a�%�A��-�X�l����b�E��(cg��[�2ֱkb��ϙ˻ނeF��.':ym�/#����:y*��`�;4z-D	>�8�,4�X�'���R����oɤ��ظܰ���4�4@&z��w&��G�+� f��Yʉq<\�Ӭh��%-~v�� 4[K5�;�=��Sp�PpXӄ,�������E0;�p ����4��C0�9���a��xf�Y�w�w������ytQ�FЊ��''!�ȝ �����w,�,-�'ƈY�6����4�Z؀���Qe�i.�-`��=d�h���ZjP�^<u�m2�>U	�fX���A��9D�0�-����<��?,��~��,���U}-�2:Ƙ��lO~v�,H����x�j#L1gm��f�-��^_W��׵$I @+vlЖ�7���U��N�s��#N�D5UUV*�(&[Z�(J��݈ˣG�Ў�i�J� <,cav!�0:�WcE��h�"�M�@��Z��q��o�2��Kq��Ld0���Ӡ ���d=�<�%���4���w�٦ۘ (<a��� �"囎Z��B��ђ��w���m�]qnUn����� <�a��v\	�@#w��eu��"��@Ò���\<�$
\���
l��`����� x� ��b��2�.�z��@PF�l��y��|2_��w��g�Z�����=6�p�}�DyM<q��g\��yoخ�%�b<�_�'=��`��a�j�.ǉ��th�WT��M�v>03�ʀb�Ҝ�'�D�x�&v}���k]�N�[�P�<����>x�шڰnu��Z��+#H�"n�y5����@yq���utK�[q~�^;3�X��)Ɣ�rQ�u�:�K�Xj"��
)#chƄ���6Ť���!�6�,&MA��T�F�̙cM���Y#��Yj Յ�s����ڇ�.X!�������҆�-����@����*�V!9n�O y@x�&t;	۔�!��}��X�P��Z�E��?	���@�:�u^� �:�3����XV����T�A��" %��	ʈ� ^fY���;�#Dod	�`v�; 5�}�g�i���h
�<�!N�|]�6��瑦�����N�" �"��B����.��K��w������~u�]�|u��E �-T�s4����.xTe�#�M�+	Nm4��9qq�X[te��f�`7f0�YeU]�E�2Y��;i����}�����x��<q�f��vO��\DH"���a��ʉ<���h4��|\����gϜ]�Dd�[4Vd��j����|@�=̭��ʾ�x���}�=�D�Y�2b�Wx�`�>=0�p -�\�&���Gt�*�İ〶����[E���R0���C���H� û�a\�
 ����^�{�-F��3�Z���� ��:s�x���U>����ahpO%�'��D6��#ܫ�闘�e�w8P$KCèwQ���E<����>3H��+���>��0 cBq����,�t��i������-b�pCݬ�h�1 �4��;E{�[5�YN�<��˴;��N�Èw����sZh�,L|87��N��CM�M�-t � |��'w����Ck<`	�b`����4}����@ؖ��v�/.x�3�:bhfnR��Cx�C�DD0��j�e�Z˼�nn��5
�A��]�J�.�`��&Q�H����SW2�1���j�]�ҁk5Ż$8��0�����Osۉ�H����}2�p �mL�>�L��f���;Q���?	��Pd3�I�m�UF���9F�0Y�'g;簘�Am�����$�A��T�����y�ip"��$�yKW+tux��.up�nL:�e�muĵ��Vɽh_�'��'ߣɃ�S�����En����I_x�~��|/�	� ��H�vߞkS)W\Ky�;r��t�Ϳ�G��t�<�.���SM%��~�ԗS͖#�:Z�:D0[�����w����9Y�շ�b
�b��x�4��c{!�C���i-�tcz�
�fH�[&^*���.���0:U%��*�LIv���]g\�^\A���a�u�E2e�`�\��߶�.�z��a��bXK�����g�@AvZ�!�,|Ψ�|�o<��e� ���e�rT��\�����ߝ'<�y.W���3���5`�n�*5.�ch� ��j�b�"ѦAV��&��"0�K&%� Q,jP�L�����YޮR��� <�ԉ��5g��q��}P]<�
��թkv-����輊���b�ӯ@8d��/Y\�	������X�7E�}�.$b�)�O��<�Ԝ�w4�>r��*��y=��>���1��b��G�^(UW��T%��"2��攅�u�<)T�1����%z����ˣJ�T�/ZO���U*$�V*��cwRe�ō�KZ� U-P����i)"��˴�b�H�`�V- �.D�)C�GD��
��!�[1C-�U�*����H�l��9�R:�b�#��ɰ<Ie�ٍ�]Q⁊�A�ʱv�cv���\�T�]tu*��B`���j��4�c9ׅ�:�-	���!0�+���S�1"�K\;����]��tή�ڹ�1e��k�U�9�X�֕�LJ�FGf��,�X-Su��V',��(�9��[��*Q0�؄K0i�+n�p�5m68V�ޙל��5`j��-�����̺���wQ���X	pl`B��[��%0�!1�<]2�3F"S4�*`cl�� �Չ+.KX]��"���rB�K�)K������D�b;v2��iip�Xu� �gEƓ֟���@A�f�G��isl�둵��4[S	#LM:ek����Ƙ�{xG���"D�ȫ��
���S��%�����  ����Ou I&�ف�q�d���i I���9����� Y�ku��c���i�H
&�t ��2��g��9��:ʕ���3І��sTR�WŨ�ce���:��l�5��O����,�z.#PXf�c�ET=�n�g, gUB� �-�p�:���
_bO���{�O�bL��Fk2[nUTI�OYk��#��"[�Q�k>a���m #cY[8��iW�rò�$���I#l^Ǽ��3�U��=��o
C��!�m�A�"�	˹��`��`��Q�'�Am�g�7�Xv2���� ou���(�_8�,rKm�I���L�h��ܢ"!$�D&���_�3�||�V��Ox���N��I�,mA	V@5�����G6�A���3\�GYY6r`����Y�ᷭ��/Cjk�U�n�t��Ye�U�d�3gQ���O�u��@��M��S��50�T2oA[�xѲ�l��]F@h ��I�;WZ�����p�_���1�(Ъ����C���yƃ @�+A2��t�;��gk�4*�Yu�(������n�1���=q-�U���c����@������ rU�:\��w��9��L�E(���Bl*�]U9���Ϟ��y���yk0[Ƙ˷�yڀ�0i����8wn�*���!i˰�:d�*���r�M�,�s<���x�Xi�� �S"b��m��F�Ͳ7�}�z�oU��o��ZY-$g	�t����7��f��T�q>��2#^�ܩS,�+����L�ƕƋ/n���1�4V��.͢��_��,�9
�?����[c��|�vOA� �-clu���[H��4�S��-Ͱ��3�\�[Ͼ�K ���A~N��{��gov" DD4@FB�e��� �Wx�������31�KJ��# 4a�$8��RE��Ns�=�x�c��Q��&D��bb�n�r����HԆ�h	������E��w9��m�q��ZI�����Q�vT1�d�U	�
����!˧]��!ŷ7
!�n��	�1�rB|�k�^*��U����ܙ�74 d���.�"�7��Ȗ���̋�g��
�����gN
@i����!��9��2�*��ekr�KEo���0{g��0�z�����`�oK��zՀ�I�u���:�\qB���dY��O�o�ME獪�&�z�$§{�Q�V�}T���^�Ŝ�z̙�3Sv��O�/�*J�U�/2r��虩uQ��/b��)�/Me�$��YPeVM]�c��o��+TZ��|2��w&�3��+��1L��r�.��J<=���_����ڹ�8Ñ�:;��YƵı"��܈]�pGw(Q�#�V�)�����K�(����%��>f uW�I�1Ϲ�s�W1w���%�q6�.��[i������|�$le�o��KIh�x���� ZR�E��sX���ĕè5�W������1�Z�O��'�l���e%PG�;É���)�ծ��<)�H|I���(�Ds��!��m���hly�{�wrq�K�9��k�K�4!@�"""O��	!ύ��aW�t�N\ A�����e�d�\3$͔;SV���� MŚ4�`UX�mB�q�y������]��;�B� Ƙ�����5[�2�̖њ��G�0-��T[F��yơgNK ,�k���3k`�`�ȑ�@Q`�v��E�O���7=츐7��8�	mo�ԫ˕=R5�31 x�c���n�4�s6`Z�󥤍4ņ�cn�K.jv�gw�P0ʎZŮ��֑;���圕��N�N�pz,<Z��0Vs�o���|�;�]d�%�n�<��>ll����ӌh�j#�;F2p�D�.�F�&��yEO>�^y����{�~H'��3����7!P,2��H=<�gM��@}��L=���1�x���t�dh��1�� P2^�w��L3#�]��݆��xڱ����\Hp����]<���s��d	x��65A C��x�C����8���r��� �D!.�&��'��G%)����DR�Qqt�Z��-̼��Fs٦m���]ca�7,Sr�$R�E�c��Vei��曯[��+M�x������[�0.ٽ��́I���]ň���O-m�(������aeE���[��p�<C`��̸�]	��e��k!�лs�{����i���,�qJ�>G�!,�oLA�<O�H[�3�> c� �Ѷ�Ŗ|h�� �R��X�����G3-<�&V��.��u�����c��N&]]x�f�8�����]R�k�bS����~W9n=%���EOKx�>c�8�q �'����L�|z������U�\a\M���a��,�F�* ��|�<F1��07K��:a�	u��s)-�{�5>����΃��j[��{קx�-�	=����׫���J����nr�<���
 � �I��0�o���4V�)� KnMe�i�����F?q�Ā,K/1���Ws�D9� %�Emʗ�"Yi{w( �D� 
]�ƨ	Ƅ	��0�\p� j��bYT�L�;�wy�>�~�O�s7]��B�:q�+M���^35�y/Jg:�xYz���n�w�4��j`�ջ�0�b�{ҥ�}N��];Pg��bLY��ƾyc��ʉ�����uYc$;�>c��G��&����+*���#&`C�S��
nR�.�W��tk"�6�J������a3��b_��8�(g'��gv�qyRIs�;W���m�H�Q  @�dM2K��#����U8�^���J�,�kV6`�Em�Sh�-��qX5�h�m,����.Չ3� �Q�l�ؒ�-4,c�M�t��4��kհ\�P-r�b�K�)a�Q�Y�rˋ��m���Q�4�-���|�R��᰽�6��l1v�ict�����-�Rh�k��6��rG&-����2ě�8�Ƀ@t��fl�V�Z�\Ce3��KMM�1�X6�2;;3R]������`H� H��z��D�z��HN t��$BO��7m��I�EPg{��q/�D*Jv��ؓ[��ؼ�m�2������4*^��5b`�@ssm�J�ø1�^q��i�c*)��˙t0����!����5����4�c�@����\�H`��Gs�D��|k�@O��������p��W sA�T�X��p�e̸]��Y9=s���n�;N����͘�ܛ��kb���U�<�5�L.�v�-�d�!�y���M�(���!0$�>8��h:�L�^��ɽ��q��Z���*����)��a��!{c����z�,���s�eC���b����(��τ�e�-�`=݊u�52a�h���<��^w���cAɁ��mn�����:��;y�H�
������Z�T��1��a��zyNa�b�<���lDύ	~�b���z�W^��ۼ�gDD�dy�ߋaݑ<+UT'�w%��Q�P�x�����G����_��wcO%�<�a�6Ž��W��ۓI��u���~7�=���.�y���J�@,h�C1]w�w��/.��'^;Ft����Į��
F�� �D:Y��J���R�)�M�nì�ؒ�0�5����1����i2ڢ;�d;�f6�Ǜ�8c,0��Z�eNO�'+ydI��]n0Si�Y3�%�l�+_�	�P�/#��~�Ш�>�onr��Xgv��01��b@�xxw�t� � �L(�z�M��-�/����H�̾>zg��^w5`;{�@^.��|\x�0�:o[y�l-~^��9�Q���d�^�j�����Z�r���� ��z��]�rZD�����/-���Nnz�s��9��h2z���ܓ�4�@�2��`�[��I�@�;����9��6��ەS������+��]�^�f�z��U�Uû��n��lo⏮��`�\x٧��^�������<#$�2%�B%��$�;åX�w��mj�z�0���Ȅ���SLo�==��m���w�|瞳�>s�������]�B � 
L��o�fk�vs�<��o��/Y�9뾯��aRZZ�%�u�6�J��)�vs4V-j0Ķ��P͖4�C�
��Ap��J�[*�0V� '�
!��6�������Ć�ܫ�J�5����x�󰰋yXpc6�}�j�h�ܮ"#��<ʄ�".ĭ�r;��zo��y��/v��7���������9����� ¾��=�m�y���ZBv�m��a�`����r��5�2�&D���<'A��$�1�1D�����	�[N������ 0Z;�bؑC�5��R%���fz�g����A#hR�~�����i���O�ފ7e]*h|V-Z�g���C,�G�su{�ڈ�7���&Ǟi�"�>���)��'���5oM���5�(E������p�r���	19j+)�<�+�{���J>QUk�yUG�"�_f��Tn��Uh�T�T�ɧJrI;��H$��&�`B@�"A,	h]r8�A���ɝm]�M��]7��qE�4s��I�))"4�2S&d�Le)�S$��L,͔��jR͚i�͓Y��34l��M4�f��̙M�fi��JnssK)��f�*iI���Y(˜ی�%�ns��i�L�h�l�j*+q�v���k�|�$��˟`���R�_R^q�-��Hc&ena��t�l6y�ڮ^�0m��A���Q{V�h�A=i�U��Der.����x_2ȹ9�(��~~�M z;�{@`Po�_~���M���Ƹ�j)nf���nA���2��̀!z�p$B��k���o=��������� X�O�9�/��{�T5`@C3M�O()w��������M�3WU�Z��R�*0���1e��l��st݆1 :̎�,H@8�ͷ+�J
<cȯ����D�Me���ޮ�� 1$�[�,5�����j�:����ވ�힇�a�@X� 0�J�X��}1��:31S3
 �r�x0�"!�
�;-c[ j}z��ss�"K�9CV��J�φ�j�U��2�@�z�V`�`s�E�����ï�/N3>��m��0�$�*O�,/3C[Y���:��T���3<�|����4�<L+�v�xP�o�zבx+�n;��ȯxz�U�[Ň�lð� M���sXoI�����ș`LD$b�/!�F$��on3	�!�:��5�$2�=��n:6l3m��]@ja�luA�q��b�;)m�����P�tA�Oj�3O�$z��T�0�8�.n�V�J�����꫟<�E��w�t5�X�\�{�����뗝I9��>�K��1	�q8"���ܜC.d�)QBf|�Ww�^������
�(��c1�����G	*��-H�Ԅtȑ��*=��1�	Qc���f�sa3�l��tgI.0at�e�����zw��O~�'��u)��f@; �P!|~�;�aաj���O�0�M��v�����8E����y��r�u֗)>����H����:(�R���LF�:&�;�d��K�f�	��\tS�7nze�Y���<L.�^���w�@8 ���c�.�en�F�w�G�h´zr�+�ᵼA�����D[�{��u�u�u�ע��{<�l���n�qU�:��U���mt���'�B q�VP[rfȊ�w��<��ߗ����֦vZO~v�ެ����cn��B	Vi�x�m��^�j���K�T�iȷ������S3-!�w.��;���H�����6I��5���vn���z���޷���s
o8aY�J�^9����r������ĩ��6��r*�Ǯk���  ��e5!$�p���~D���|�dm4qd�;׿�������iļ��$dϲQ�@������le�^�˟O-��	c�bH�\�H��b*BU�&�&�$*�EX��!y�\渺�5S��&�C�*���D7RquiD��ݒI��F�Ze��n�Z$��"��f섑�/D����	�AL������*HF�i$MYRB95ZH�F�K]s�mhъ��\\��[Y4�� �5SM�f��G���R�κ�C�k���	:�qS�����Q�4���`9�w������{g+IZ��-kmE��+Z�M��b�? �~I�"?_���~���;�dplo�܎4����3S��xk�x5���K=�mg񜸞�)5?�9x����{�����q�=)����8���ږ&�P����no�y*�i��=������i��:O���i��߷���s�Ѯ猄=�Z?z5��:<��T�?���cÆ�����BuG��*!"G�F�E���I�$�����;<�͸�����p}g�=$�!��蓏�L����f���Y͞���>�.㯙���|��S�vW�_�"[�!.-��S�}NO����>S�U���x�莴s�G�I�ӧ������FO+��.,�%ޥ��lO�X����v����d��#R#��r7����'N|��0�O�k��jv=��i�p���ǮG��/�mn�N�z7~��oZ��ǻ��9����[����h�kI��q$D*RKJ	4���Z�Μ��(�U���%k\��\������[��ŬTj6�KJ�ej��XY-��,�)-�-��d�U
!%J@�EKTmF����-f��m[M��i�mj͚�M�k,���m��6YlY6M���E�fi�-\�3i�4�IT-H8(j�����CR$���Ii"iQ����R¥D�:D�ҵ˳N�\�M8������;�u���7�u<�:���o/�x��А"bj�����x}���z�Q������I;G�5����>hL��VWu������z���?�֪�-xC���{��O$z����܇_�����=Ge}i��^���������#�I'��M��h�",h��ƍ4j�ѢƋ4XѦcF�64h��hƍ4X�bƍ�E�*,X�b6l��Q���ƍ��ƙd�h��F��fYf��,TXѢ4h��ɣE�6�,lXѢƍ���3E�,h�)�E�4m3cF�4��4�,h�*Ke�F�4�ii���ƍ4X�6liJƍ4�Dh�b�Ѧh�4�#Id���Ѣƍ�E���X�cF�4X�d�bɤ���QcIcL�cF�4i�Ƌ6*4h�4lh�cF�j4X�bƍ�(�cQ�ō-#F�,h�cF�4X�Qh�cF�Ѣ�cd�h��F4i*4XѤ��b4m&����4Z4i�L�h��Ƌ4�"�54XѢ�h��*�ō4Xѣ&���4h����F��SE��bf�4lh���ĳF�,lh���4Xب��ccDh�bō%�%�F�MM,h�H�&�&��F�4S4�,h���ƓDh�,h�ѢƒĚ4X�flZ,�4I�E��ƒœE���,�,h�cF�4i,i,hѱ�D�Fʚ6��رcDi�,i,Y,�M1�bƋ,l�M��,i,�6,h�4X�cE����i�K3EF�4h�cE�K*4i"Ƌ,h�cb�h�cI��FƓDli,h��řcD�4Y66M*4i$����ƍ%�#F�,�,�,Dh�,Y,h�cd�,lY�4X��b6e�664Y4i#I�ƒœE�"ƙ��ƍ4���cIcFō#I�Ƌ,�,�"ƍd�lh�X�b4i*,Y6�4Yd��3E�e�$�K664X�hѢō*f�,Q�E�EF�Rc)1D!Q��2`�1i �2%QIF,-�ѱ�J�|K��e{~�5e�$���
�2W4��8�8|���~c�{^z�kT�����?'y�W�ã�N�s}y!���u�����<���GI׌���=�I����W�K#�o�����L|�������Y:����=ozH�A�⛲|iR��Q5�=�_t{�[�r��ϕ��u��CN��wu�v��W?�*(��o�>�䜣�^:����´�/�z����XiK�_r^#Z�OK�$�O�܆O��J��ގ�4~�|l�h�!�-$��9I9Z|����-�R�<ȶ-�������#��$6�q�8<u$�H����uChW(�������D���>x�'�szXY̍��:�:G�M|���Ԟ�;��aދ�fڅ�M3~}�  �a����[���z�'j�e�;U�$�R8֤i��w�j�O��uD]vO�'�>��$I �����'�/�<�O���R��'Æ�<��'��>����?tt���s<���О����88�T�#d���|ޯg��4,z>UIc�|bt�Yc�H����N��!������|���d~��4�$�voey�s���KV�~P7dU��>��4���h�'��#H}m�I�3�i�����N|��'�������F�O�:#�JK��)8�|}:��?ݬ��U�����Z�w�em�_i�}5<�t>$�N^��r�wf����)i(��ې��"q|k��r杵���c�p�7um���#<�6w<�o�s��$�jK�}�oZ��X��4�5�zռ:Nk�z^���79NG��N�(p�RQ�v9U��y޽]�rN�N��گy��w]iэ�잓���rG��ďD�eUvw翽��wO�/|}V*��#��o�����	$'�4����'z>�h��Ji_��8��|��睐�B{WҞ��'�ꌎ'�N�>H�#q8�W'T�X������u>���g��M�^�?7������L�D��c^<���m,�$VI��/ZG�?�.�p�!>�3v