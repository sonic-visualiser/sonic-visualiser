BZh91AY&SY_cf|	�߀ryg����������`�~    (    tp=      p  v;}
 ����E(P� 8Djͫ5��	���8�/9�h���u΍�.W��4 ��X�)��4h�:(2ˊ::��(���qB�<.��7.�(��C�G�U�s�(��j��l��]oN x�{�g(P:�\Q"�8�Дͮ(��qES�˔P�E<ޜ�
f����CB��s^(Ѡ9�qN��2�� ޏL�\��V��(���                 �  P d�T��L�4ɦ� @ɠh�&M��R#*��#ja0&��4a40��i���RDʔ	���� 0� b  )�TP�PƂ2h� ��4Ɉ�� A
� @#L��4ɦ�M�z�I�jyOO"G�j�~��&@        ���C�<_W���DBO��8���!�'�HW�� �ވ"!�tU���������!�x
��{���L����|y��ƿOn3���C9�������'��~�����������Ӗ�H���Ⱦ����N�D5�ێ��.h*��@�B�iUQ�bT�&1U�t����ǧ\2 �>wU9m�m������zk�;��Yɢ=d�xc�錝Ц �Ӗ_�'�;{:Q��ax��֐�� �;p��(ny`���G��}?jc�����|0n��:��+�� o�>c��m��+�������?_ٻ���-p$'�Uw��{�8�H.'x��(.�
�u	�P�!8�P���⫡\	Ą�Z�*����sx���N$
W`�H(+p+�8�S"]	��(.

����{H(.�'�	���p;���H.$

�
� �w�W1! �
�2���AC���N	WBBq!!��'�����x��HU]�Ą��(.*�U�	Ą���'AL���PP� ��P\<�HN$<d8��N'��>!�A8��HHN$$8s�W{�ؐ�HU�U�$$8�W|	Ą�BBq!W�-T�	�p$��P��<�nWq ����*��q��	!8���\(x\�U�$
�AITí�M��lPP%�H.
	p<d/*�`���Ą�BA��!!���
�	!8�PV�UPN$'
���]�����{����x�	4!!8��n(7>+�=!�Ǥ=!8��!<C�C�
�Ă���u���
�$�&���	Wq$�2��v�� ��bC���q8�n��]�{ۨu���		Ą\	��	ćk�H(.$$*��
�C�9����HI�'������p*��8��U	Ă8���BqǕ�U]��	��BA�8�\(N$ć�C��z��q!UF���m�=z�=8��!ǈHN$'�p'
�
�	�B�Ą\�q8��N"�N'd$'�HN'��	ćD���(H5w���p'�����7�Oaa����N$$'	p'!!8���BBR�H.$'��"�!8�bL�!	�$%��HN$$'���		�!8��	�Y�^�q8���C�	P�$���H.+��D:ܼ	��BM\Ą�BC���HN!		Ą��p<AHN$$'㌄��N$�N$!���HN!BqHO����z���$$���HB! �1N*��		p��{p!Ą�����7�	�P�b.��BC�<��9p'
����p'�|���8�����Rf��w%�   �N\��M`�u�~:�}=3����O-�����/O��js|M���ז��xq���~���N�/�������0b��@�[��l��r��d�D�N�h����݄�@A8,���� �&my����FiS��L�Ur���b��/RqŽ;�\�[��!�Z�������q�p:��(�ND�QhX�i�bLC�A�y\��6.TA�xi�q�8�a��a���Lࡈ%# �Ub�!H���s�6mN5<'ė��^��P��;�t�bk ��~J��:��3"&L�\�hG��R�=>��d���7�P�0��OE�5�@��h�=8%��B��s"c��$�R-��"/�ż�SǢ�J_��A8���Xj�'� c���Vn�PS�N������uF���t�"�T�UA�X��U,x�T��H��4�#Bn�74��}���yf�ݥJ�.��I>�(��MML�S����p�"�J��#M�8��Bļ�u�9��(c+#.2br��̡�����Zd���j&���{Ö]H�"&&C�s�nd)�y�up�Fh'jOt��3SJB���C�.�7sx��[��ZyF>n����GԽ�w����j��.g%�1j5FiM`W�N�&2�K���62Մ�O6T]�uss"q�=ӽ,� FL��J^��6mɃC.���B�`�dEVfd�e �j�vr.
S�#$9T-F:c�)��{��W�]�jt����SBdŽ���������j�(�@R�W�Ō����x��P��S�r�`�y�zx̬���
ѻ����F-�|�Of0�A�� �,�H��_�7�%]܈{|�b�&���ʇQu99b�*�Tr骎V9|k�_.N#Vb��hL��Z�{Q�����)�&��P%^Y���c��eA	B�RN��e�FELe��3)�fDI� ������Ҫ�os�5��1�A�Yk*bf{�*��4.���\�е��I�DJ���#2�Z��ȻN��"�z��$��#�x�/�
��u9�2I��S[̫��汌�.PD���qs��d�&����Pt�L�ǜ�ȣ�L�=�������<(��&.\D���PI�LT�<���Q�[�W��'�Č��1n���+1LTeT@���ɀ�	�$a�w���\K�L�UI���H3J)F�/*o*��-�]T�W1n_�:����rl��X�Xr*�Iȋ�wb��f:�d�c�������UJn���.�>H����#,��T\<*�!U��0&�Ud���D��
Q��,]�	�J����L�S�2_.�o�^����#�Y(�D��2��1/�������B�ٴ2�\�Ž̧�D��FUS��nս����Ԙ�sbMM̄`��B���(�����9Riࠞ�T)Y1Q�tb�����n��aM�)M�	��Z˙w�D�F=ILd	�&�JyS��7	�V�Y�ǥR^`**-��(RF������%UW���e�.�Ip�3�9���eD�����Ne�ɁE�Rqr"�ɑV&��*�����p��y	���˘���o"b\�Aw�{�Tړ7Ouu�%�.�|���P���$�S�	����^�E��&f/؃8��z����4��!A`�w|�5���WT)�c�`��0���
�b��<�x�ÈM���R���>�d�lk����w��O3�V�7T%���*�0�J�  �`� S.�6e��&J	v��  �+u� V��	rX �HU܀
�7@�` �X*  �%�J�@eeLA��
�.�p))  $D���b�Xبa�D�ܕ6�PKD7wkD$Z`K�Y4@� "�]���
I X�Ar�������
a[��	��I� � ������(,���H6f�!7wK�A{���2�!��*@�AHU�@��W.��+r�N ������&��������5��m��%ƕ�ϣ����&/������GW�@�; ��ˏa˗��ÿ�g��l��xp6�9�'q�㙵7��[�~��B���;3�T:&�x�O�,d!!Č(S�6	T�ۺ�$���?c�R~���^�h|9^&Ƥ���m�]�̻
AJH�����Č�����o
1q�������aHUm�-� m��"#`���Щ)��B2�و�d�Z��B�Tj`�\�MJ�G�"�c\]-G�gR��E�wݑ���E��h��fS��R�3Cjnc#�kG$�Jp��A6�R�1�矷��]ې�T+bY]4�� �������bjYw0MT�ѷ<(�jd*j�R7%3[��1�6,��M�MSv�������U���uó�9��ηR^m��k���P0YEK����q�j�F���	��cfUQ��.�4�Ƙ1�.���6tJ�a�3H��b�\:��#ܘV�Y�������DMkJX#@�R:�T%�v�r6�R����]kM�j��\�.���������5!��4��K�-D���[��b���L2���&-�U�.�j�h�èdhW�q���Y4Ta64��ghm�]j[��f�/1���b�6�t҈0�jL�����U��mu��3+�Y�	��u͸�Z�)C%���f�hU��*��6�Dvlv�ER'�ݷ�/G�6ѫ�K�hU�� kMdõ�J�[%� ��[Q)	��(n���b�j����Cm��%ݺ����@fFg+!5��Фt���9��I(J��3�ą�gMK���6�-���m2������٬�h�BH������l����b.�!�D������z�[�X�b���Z哴?zy��TT���`�h�"W6�CV��l،�q��r,3�U�fֲ^̲4���J��-�,p\�b��Ғ�yqv�4&���gW��Ԕ���Gi�5�d���`�J����]1V�$�)m �Cs%�
����;4�[5�e�ㄡ�0��4�bXk���8�WH��i#�5�`��7�v��b��1��X �mtr�L4n�qs���ZS\V���J8�+�GZ����h�Vm���- �R�I�#��4���)E�\�l�CdB��a�S��J�����Fպ\�15��掠�\3Z�h	v�6t�+,js�o[Zv�m�z9�l2���B�4Ft6ؚ<����-�$&KMur��^}X5�����{��k�pt:q��  ��4���nq������"":��u,q���:m��T����NC���ߋ�G����G'|XN��_��{��G�N]/w��_��yc�0=��z��m��T�0��at�����3�DZ�Rþa����$���I������EHN�@���X�� i˞G�o({ᩙe�r�!�y�t��N�GN=ս���������=���{i^�Ҳ6�G�RI� ��4����:q��|^��E_R=Ȭ`XD�$�Ίy-�y�GN���өa�s	ڳ��	��y��zi^�%�^F3��B4�۽�ɓ�=��\��A���ޗ�V�R$aU39��D��t�'�xS��~q==�}kQ|=n�_�x1�;�4���#1+}�M*��=x�%�S_|�<�Є�5��wq�\��Ms-��ޞ��z��Sk�!�&�g}u��om�Co����z�y�}#�i��JѝN���ȁjL�4MS�A��$�Qi(s&�Ϡ@���]"H�(?�ǋ�u�V��d#S"��sI��\H���^�-)�8(ZB�&��2��Y��U3p�0̄����w��~Uzfo}��e.}��7||c.�$|���4����,���SKS�Nݷ�������1:MÔ�22�8F��ȗ� ∇�
�o>�8|�<y2�����c��e���_ϙ��I��*��qFKdӹ�aX�����n��|�{������m��%�t��&r�Q-�B�^E>f�FH�b����Ԭk��[��N��wm/��=�T��=3u����O^���ׅv��t�*��Ř$b����=8�G����i��s-�}L�c�!d���y	��E������XR�/v���y$J�U�[�!$k<��ϫ��Q}���kI��Y���������mv�t��.%����go���]zI�kf�s-��Q&Hњ�cv��J['�OEfL=	]8V��ޜ[���{���n,��G�l�m���>S�K�{ޝ�䁝��a9
�D�g#8E�y�qX��K`'�����{�+���x�Gn8���J���c|�����\��bD�8Ը1�4��p}<O�N��Ǔ� |Hz�Ï<�/Dgt4�{�N'G���g��]@�$��>o���a���{��d>����g����t��^�<w�w�w*y��>�^��q������d��=O��CǼ��g��Fh[	�}hgY�C[��3���=�p�|P<�P $d ���]>L'��#��*~O���吪(�f�e�4 ��E��Z]��E�B �0R�7AH�  �L2 �(&�*5`�:��$�]����ڄ�����~��Ņa�6�`ܡH
��,j j��W(�T@P
YM&�� lٲ�� .���Ү�IQ�b����.�Y�pd~�0riޡyBBͪF����E�;Z5�҂5��wFw��.���ʶ�Բ6��L�ٚJI���ZL��Yn4в���$+���ձ�m,�
ji��YXQX4U��m"�k[��m�+7g6fI#��J�X�ґs�VE�`����Ep�\Ĺg�f�L�Q��@����3mpm�
�A[CJ�)�F,��Jƚ�vY�j��q5�V9���˴���Q-�h��M,�q6�p`,�O������6�J̊ҍ�"R�a\IN$З0Թ�b���@���D��l҇���'){US��*�@�(![�f����Vq{���r��!M]*�r͎r��ӱλ#���ᅹm��0�i5p2S�f�f��1`H�d^�:i����G������V%��X���+��� ~�K�a|�n��2���*����@y��g�i����z>�-�K~s�翞�v���;�˶ÅjA�X��x\=;�`= qf�OQ�|h�	ϊ��Q0�3D��O�M���s�#W�gjf�[N�l0���V�������7&Q�\��i�&�O��a���00���@����׷��4rEP��qfH%��R��o-�X�&vY���m�	��z���S�cU�:��Q�p����z��R�[m^�`g�W���V"O�k�a��8��z���1vM�E�5�n�Kc]`a��-��L	�!(tRQ��:O����m��1ݥ�K
m v
�{���7������8M�'���ʝwS~��>��\ P����J=�u�18����B�^�^W��*�6nf"�5M�nWqt#.��`M/�y���(�%d�����V��`c+W�'��c�n��w�JE%���(�.�v��ʶ�7���>�oS�ֻ50���;��+m��:�޾ϵ]��������&��.'*I!����Cz���F������4	����"�٨��l���!�ݿ9 ����}��l�ߜ���;_R^���;Lk�s���u��f�N�B��0�K;����j�D��/�뱗��Mv�h���a���{n�z��^C��6��fD��ۑ�fDpY��6���I�9�Ml;z�G����_�Lަ-��p)����m/5�/kь���@�D����Y�ճP��<ʅ]�"� ��rR��Z#��n�z;m[Noz���zZ�
�A,k^U0���}ϵ;���N�y絼�| jĘaH�	l��K�	ؼ�6jw�T3	!���א+�5$����?�9�`�[��
���%��u	t��yO'�*�"��dH�%6�@�;i6�n� &�0p�l�jF.@0V,����O�7��	���kf4��r�4��lS6߄�^U7�������յ������L�{8&T3��ɵ�����x1:i�ه��T1R�]O���l����:�M��M�ێ�i�6��) J 0��֪��צL[��v�7ga�ƘKm��'��l�X3<�(O�5��c��D��&��9�r�N6�G�ٓ{�n�������rq_�V���I�,��y�?��o�y���3+�$�=�fL��m܊���$V>	w�Ly��J��]W�z|"��ا�)._�y�&��L�Ņ�Ag�Ib>G�5љ�yx���ʿF`�x)�'/oرO�4J&��_}���}D߁iu�2bc���c)z�s4��?��z�4�(pD0��"�Q�F�<�(;�<9���w7�����r�uI,~ǣ?�g�a��If��\��c�X��x���1��yi

IA��	��×�a�xU���8�n�p��p5���9�J�H��e��si��6�X�b����Z	*�O *�x��=<���o�`�,�yCq����C���2� 9�t<Q�%�O+�@�1�ƕ�?r�Q-�aVt��wz�!Ő6̭ͬ��y�M��� lΖiZ���-��������z� �%� ��'�(ި��]n��]No��D!��1U��0kW�z;%�gR�j�%q+[d�b�!d2+�)%�,��a&M_���@�kf�����AVA҈xxv� � �h
���rA��E��v��8���ڰ���=�f[ �,�-Z�l���N1-��?����Ǟ�;���2)+��C�f`�4��	���ʇ�n@Ȑ�rމt��d�f�H�d��_�N�6�6dz5�M� [���4���#�x^;qE\w4���s�w�/Èw�%<*oc�p�1~f�""t�cd9�4�\HE:��GP�H���/�Ѓ���oz�2�-Ly�d�;I8��|l�y)�>b ��c�]/�p1���neWk��䟩d���v��H���G��sG���8�2@�l`;o_8 \��(�wv8�nR@��8�A�A��z2&�Y�N��B^�7n�CK`�$k����'�4[ e������f.L��/�/<�|apw��e��`el~� �e����:ZM�t�!�v�B��T���Z6s�ͿnW�;�o�'>��U�W? �A� ��w=꧓��oL����~�8뺕�����1�!�l�������y�d`���;Y1l�ºY
��|o����^Fxb���'�y�Eq���c,vCjV,nǇ�}�x��PT8��i}�)n�
��2�7��KYo�q���Q�z��-�t�U�ql�9}r��睟O��.��b)��Bw�r�ե��g@���!�@tIǸ�y����U�I��	��w	�Il�n6{����M�[�0Qa�X��y�U8E�X��`d�䝮�5Q�hf��	<��d���E����y� Z�8c�H�w��Y��=D��r�.Ӱ�)8^sݓ�5J^����:�;�zSጚ��a��Ѧ�x��3��f�2��
���4�mU�OC���>I�y<	=�2;���(�c�[�j[��,a� <־���B6�`��2��Y�h�F\\)�Ox̧���<�b��j9�4��lAJR+"DT�YW��H��w �>4}��{�(,����p;o�{�Q�x�i�	v<����L5��$J��a sh[�Y���$�a�X�(DX�Ձ Q DE��1�J�K�
 Ո���%�;�ͽ�/ws	d�w�^�fd�X�� ^bs�E\����φ]��;��ؿy����>�j���@0B>�2�")��D�M<dX����/2${(��<��Q�^�B�췘�G�µ�f�<mHw����+�;Y�������F�a�z<���S!M��X|/��3�3�L�W_/{|�|>g]\͛��z}�pHH ! 
ˢ��@B(��  ��""&IblF9V,b��!>�y;	e��<�.\:�&+�s�kp�f�2�J� v1����%��jms�mQ�D��Գw�t�Ұ���2��:0c�K�̎,R�U]��%�J�6��![e�5b�ʒ��0RS��i��lŴm"l�E��������1����2�Y���a���)5	�m���Ms�6�Z�j��l����6�)6�CЮ��WlgM��.�c9l36�kE`�%�STދ���?O_�L����&�W���}�豨"!�h�����*��ϒ�gu1�b��&�h���XX�ʻ,ȅ�1���d$�$a�M����/+.�p������w��y�7��!@����k�ij�2�`D��d2�Ø�+�'�a�-$^�: %���4��&-r��`�4��ã������κ-F�Dm媻Ϝ��!�`V\y��|�4�F�t�ȎY[x�λ��Z�I��)���D��`[6��$�|�e���0)6��6p;��*�����w���㖙��u��t�$�C�M�Q�	��u�Ĺ����0Ź��:`���RU�����,�F�h�N&5�@���ҋ,��� �Ō��v��-�Ӷ�=l;�x;��v���,3�\�rHaA@x��H	���	��Rm"�{I���$7&؎-GZ�-z	��@S7݉�/?\��w�(A�e�><�F���\\�����}���
�D̕�W��{��<�ʞ��U�{~�t��Ӑ�[����	a`-c��k^�@��8��%�I�-ű����zuU�"*P��~"�̑���2��s��U	�����<1� ����ݟ�S0�v�lh�vu]5�&I`��x�)*�I�Y��*)3��A�ʬUm�W.$�Db�"*Ȣ �egG����ӌl��<���	$ig'�4=�%�y)�T@��;�ʾ�i���!����3ݝ�{��,q��Q��P�$��.�����{�����W{8��Y�#C��ť�q2U����u��[��KXʁ$ih�7rǳ<@���b}����<�=#��V�8P�3H�X��adl�Oc��`A���d �Go=��2Ǥ�y,ʰ[��:�,?�5�`�F)�8t�G���di��mc@�;nx< �@��9Q���N�")D4�:u�67��YX� �m����*�il3�x��s`�X��Ae�g���0ܽf���A�O�ӧZ���w��nE�a�8��<@O>^Fϗ��Ɇ�s��$�,<h�`���K��5��!wC�� ̦|���fXqʾ�{u����l�� � Q24��8��pHPv��;�^_/8@���h* $����S�ίs���զt��Bh��8Z~��/��FIn$�����T�m��z�X��m���N BJb"�1a �Gx���r��Ζ� ��.�:Ũl5�"�h�YJm�QM��OM��@��Zƅ���'�g�6�{#CKVd���OHd�`C�[O�Xw�Օ\C(1��L�����b6�^n�\MjY����1��%�P��Z �I��8�F��M�%�o�32 $��FPΨ<ʧ�(iϗ��S�=|�s�y7�!� &�W><�"ZP�v;R��WU:"jD<�q	��z�ס�M�5aE_�<�竿x� �h{ ��ժ}1r^���[�4�/l	!�$�������_��N�v�Q6\97�n=jAqC^m�����Z�N<�/T��N)�eR/5�O���5h��>V��-g������Q����Br���
>��+�yA]�ӣ�jf=+=d��r��C,�p�9�������Y��B����"A���JJ��$@�Z�-"e���+p��i�|tȮ�'�Z�,h�^�5}���%6�IJ�惌T̈��e��4d��C����*}�zD{I���b�6b¢O��%��������r���Ӝ�0���,ԅ���&�-�#.m�S�3��~�m'{��P�@Z1�J�.QC�
:l�᰺̍��m �$�ѷ�[����$���AX��ܲKi-i`�g���� Db2�XQ�3��n]�Ϝ���=���6:�u�z��� ��(B}��뱻5�%V�L$GR��4�v���!:�V�$�Ac���j덓a�ɍ��g+H2�edp�l�/�O�o\�y�띧q���S�R�y���6�a�H���c�$Qm1k��"@��%if��@}ނ �B��xBt��()9�������D&p��$I]��g��<QE��w���;Jm^�]��b��'C�u���Q��H8��3�[-��H���x����%�!9�H�C��c��|���=����ګ�@�͆���8Z6��lq���&0��8Q�U4����B��1��j�k���~��n�n������mU���j��>Y�� [�OO $��d�tقӧ��y���0��lw�z���f!�(���0�ȱ���f��s�h˧ב�l��le����YǊV���snL���]��\�(��&J�q=����8[D���e��� I@x?sۉ�
:`
N�vL��9�0<95�0ޗ�"-f(��o�q+/.�sv}묜��_~w�m�eA�V V,":����-]Q�vu�Yx��ۖ�Yf�M���8��[m��Rr�Ҳb��
�c�b��\-�����~_��Ύ�{S�q�2@7F��y@�Zl�> ��`x�b��Hq�M.�-Ǝ�;�������D������w�(�qDa���u������{�T ��=v�o�O��p��>*���,�ۙ[����a64�#H�|#U�Ζ�&�/�/>�~�m�%W���!�P1� ���y�"n���L�o��� Qhh�\��	�a1C�i�5r:���{(��\=�Ӊk��C����<-��f}��	(f��&��p��/u��<���������e�m�I��P��A$L�4�s�6[N�e)a�	c��RX{�?n�Ȭȷ���h �3n���R8�7g>Y�>|�w��c��]�`��T	�y�h�p~d�cþ�@��y@�p�~?s�Ķ�GX)��[�?!$��-'L�!�;���t�T�4��Dhl����qk��f4�) �J~�9�pՄ�d���s�$B��o9�&��@��9�s���D�����s�� t�$�?�ř��r��\����tfU�z�Ԣ)� K�x��^�?�	�u"����≊4��I��
����ǐO�ב�w~s�}v�����z.�ÔdU��Z�V���EZ���y
� ��]ýқ.�[׎@�z�D��Z������=Q�#���mQSt�
q=O��������������c"Ȕ���T$��Y��
�R����SWE ZR�.HҫR�+��! S���#*��>i�^GԾ[.=$R(cf1��ݡjj�P�:݇�����tH1�9�P�,]�!i����Q� �-�J���avM�׊KV;q�\��e�]�,�HJA0�I��j�����\��V�ͬ�e����������J�h�H��YFVT֍��]0���6*��Hɩl�i&��ʭ�9uKl���h[�Q�nU8]l%x9�#���[F�nmM��w,4Ɇ*�h�s�R�ژni������^��Q@S�ؚ"S�8���hh
(b��B������JBbF��<dCY��j
���r��o._�w��H5d����Qr�m�B-��X⼫�_�3��vvX�h��"�0eJ��%�5! ^6��헤�Х���i��9�s�)ŭ�<^CRl,@���<L3CU���e�~|���i	��m� �\zØ���Qf�}�g�� �����Y���� �I[����}��vIظ�j��YTT� (����	:@`>4ZH0��"���)��O#���WL�8d6��׳>-Dq�`�m��>c <ǀ,��;o�#K3 Q�d|�O���]��0Y�l�2��y>ޱma�����n���+:Xd)�W	�:����ځq*�
�͍�0�c �z"Y�BΖ����\K�����r��ɾ����f0Q��*+���r4��3�R�y��(i���-�K>�~bH�7:�/�l��'Oa#r^�q�\t�n���C3{[-��sʿ��>����^��d��2�nj^��v���N�흳�7;]��$�X���4��r�6��Bou�`�v�� �,\���io~X�f����/eo+��L0� @��G��ы:s/�xo��'� D�LD�.(�M��˽[u��6]�W"M
g\���:�t5d"V�KJ�\A���3�x�@���i���@�Yz���)��1�
`�!�'9�r2=N��|�����n�H��7|�@r0�� �p��,t6|�y�ñ|"�B��1����q-�kX��L ���b�e�D<"�At
�N��H����V@�<�s��b��=��X��E���,A��|Z�Y� ���7��[Ll\�XZE{%��g������j2�]L5��0j����='~��|�9|���k��8�-��������H(8,i��s��_�q��ݸ�.-�r�Ry�5��8Z��!f`��(�}�`� �̈b�C�P���m���k���9���$�;Ӡw,�,-�'ƈY�6����r�w`W�N8���>f����OY#�-8�V��&׏`L��B|[�|��.�����V(���rഏ�Z��%�E|Ʌ�������GX�m�I�o����I7Us�-Di�"�,���Ű��l���  """[�f��$^]�=+�ɟ;����_6���s��V  #ou�Z�D	BW#0�h3p��&���ٹr�HJ7dq	/ᖳh��U��l��[kz����"�R���9-��o��N{�,a{�٧@ Ao<�{�y�Kqkia%6�[�M�0@Px�G�@)vE�7������1��R�LȄRI��NJ����DLL���#5���O�`��+�l�~��^'��� R�6@X-�Sd4[L4���$O���7�,��w�ϳ�}�w{�G
�AI҇N!<@�!��~�ޢXa�l��[~ ���������}0#��Ś�P�y�ʷ���b�$����8��
���}����&��ѣ�a]S�;�6!��� ϫ*��Js<���������ͭw�;Qn�C���dd���F#j���Oqk/`��",���	��b�S3s�Ǜ����/�m��1x�ύbJ�P�R��	F=׼�u�lC I%��I��j�"�h������(")iJi*"��")Z!�)X����j&$*����� �)if&)���$�0a�MI�	�*��f����-�θ\�C��p'Ź�6[�s�b� �S
�'-�)�t����q0���Hܤ���ϼ��x�kB��|�K_ ������#��Y��GX.�"���g_�|Cp��
߽�=�<�N:�͗b/��,�3,��S���7���;Y��޾�3�4��L4�x]��i>.ԛd��[��'��]yW��|��=DH���6���O�����'�g�����~w�]��w��E �,�s����.^s£.��]I08�zBG^ee��U�A!�[�1�)���m�0�A0���Qr�(��d��l�x��<q�f��;'�{�"$V�Ű�oeD�KAv4�zy>.CI�n�,�<�� �h��qF�1@Wq> I�V��e_C�<tz�q��PԢqK��1\�ݥ������L8�� oW;	�e�`��&J�q,8��y��>������{�ݪ���"���s(�G��z�a�Tt�`\{���1jcC������Ϲ�b&�T�{�=��ahpO%�'[U�b��r��X�Dy��^�p��"D�<:�u#�c�2�O<�o�ό�3����{Ͼ� ��Мp=n�'�`6|�k�$�(��X���k;!LD�2%m��^��@A}V@S��,�2��"�����'� ��֚  ���8���#M�M�-t � |��'w��6��� ��&
�q<m�0�sG���}��V 3.�%�z��Ν14�7)z�i!�r!�""ED��k.�5��jg�U��:��nt��^fM#,")��ˡ��6�A�j��j�]�ҁk5ŹCÁ��#	�L�+D�=���QZ��p���, 1���Ys��]�kɨ��D	�~��0��gF���貪�[�0r��`�TN�v�_0&;��[\��=��[o ���*�k��qŋ����	A��o�����:�Z���U7&d���6��Z�ykdDo��ϓ�яd�ލ	���ecA��9�˹M�Cy��|���� FL	���o�5����%�㝹C�:afߍX#��:N�@k�yک����ſqb(���e�~Nt�T<-g&������w����9Y��	gQ�Us(&JcH.F7�P9y�6���'F7�ప�d�5�e⬯i2��0�)�ҩ-L9PD�bK���:�"����x��2(y�/[�Z��>���K�ޢe�c0������q��g�@AvZ�!�,|Ψ�|�o<��e� ���e�rT��\��Vg��;N���\�/��g��ҍXa[���K�DX� j�!cZ���@��i�Dլh�� DE�&RɉpK�6� m�|�����޽�m�߈�ί�˳�՟c]�[��At�H*�V��Uط�/[Ӣ�*����N� ᒂ��dQs$&8Nz'�^��c�]������<��>���Rr�����dL|t�n��H�����^��R����A�x�U^��P�"�ˣ�R��X�S ǋ�>����W.�*�S̽i>Vb�T���X�lk��ﺓ.F,lZZ� ��j����VHiH	L&]��2D����h����p
1V5�EP>����æ�+ǔ�f�l��cYWP���۵#��2��MH�������&��%��f6muG�+)[.�e���aH`���Zk�dX]q5l�b(�k�l%�YXμ,��XhM��	�(f�R&�����l����SAvw u�:�#�j�lŔ3f)�3nm���$��$L�;7&ҍ3 ͨ��%��nӫ�y����al�T�au��`�6V�L�n�d�Mt&�￩�x18��z��H���"�~o���M���!���s5y-�bS��(Ɇ�n/Q��œ%I���3L`�V$���eJ�"��dsP�荳���=9ܱ��1���rc)�N�.S�k�!������z���h:l����­.m� Sr6����ja$i�i�L�~yԻx��o���ggcv\��[]p��i�8*�c̤�o ��n'��$�F����2	S�����$���y��Kp��k�|���]n%X�f�ZdR��; 71�L���ݔ �����"!(@�wwx.����Q�<��p7�u����k��A7o�Y��\F����Ǧ��{B���.X@Ϊ�<�L[��-�uO)n>���3mp�(�	B(�u v�f����>s|<�~�Ͽ}+��|ZϘy���H��؁�u�;J�;��Y%gH�
H��b�;u��f����=��o
C��!�m�A�"��GV�+[l2�'~�6O�7��Ϗ,;	:@P{���``��!Gt�*�āc�X8�n�L��p'����g���޳�p	 �D Z��A�zpK9jOd�!��""���dn�&SV���c����L[]�b䆑s��9t#��e�i:N�����rr\�,���L�l�@$�J �fXi�x�D&�m�����Ū7��	��<h�m6dv�� 4 |� ����HӾ�g ��
Qܪ�Gcl�6�N��|���Y;˴+�gO�	� z��q���}�}�3�29���9�l"���Ņ��j��-gKA�-:@䫞t�%�﫣����{vQ+0�&¬e�S��������m�<��-�Le�ۼ�@s4��@;�A[V搴��hi�\���˩7������1�Sia��߳ߑ���gU[�a��h�YvH3\@���˱��C6��ZH� ���KQ�-E�o��́��X��"�Ȍ	{�r�L�0l�S�}2W<ߟ>}�=� w�c\h�@f]�^"�� kB���ik��ǣ��0��gŀ>X�m먖�(��F=y�9_n����ϕrmo^�45,�ff�r���.y��������<L0X�W�����"�F��bS��e6�ѳ�֪�HF*BQWE�"<�glT$���7��cln�sk�#��\;�~R�{�_s����ߔjCM���[��Ţ�m;���]�6Ÿ���$��y��M�(��*�6<��p7+�*S� Rz��'�y��7z݄��9!>w5�o�*�yz��3Aր�;�%ײ.Cxѱɬ�oo=<ȿp��-��o��N@|�]��>��/=�@�aqJʲ��!	x�4�%��=��hս
G{��勰\7���j�m>
�����O�d���B���dY��O�o�ME獪�&�z�$§{�Q�V�}T���^�Ŝ�z̙�3Sv��O�/�*J�U�/2r��虩uQ��/b��)�/Me�$��YPeVM]�c��o��+TZ��|2��w&�3��+��1L��r�.��J<=���_����ڹ�8Ñ�;eu�����%� 18YA$B���T��poA�1���on{<7�]�G�Oq-�Q�1��hB+�5S5FܵDs-[U�Zw�|��d7_\)���H��n�;N��4�h���Bjt�[��co��W��a\�Tkއ H�e"�w�T� DUvL2��#ˁ'~V�ݝ����[X��>��|�g�t�"	9����6�Hh�4F��> N P�]}����" ��ﵲ������󯗝��}f}�'��DUW-ƈ��ڜ�p̓(ۥ�69�]�wRǢ�a! �T�[t�m��,P(G�̷�(�M�L�5�: ��䜾1�9Y5[�2�̖њ��G�0-��T[F��yơgNK ,�k���3k`�`�ȑ ���w�xx���Hu@i}��χv\H�k�k�����U�ʞ����<]����ͷX�x��	�0��~y��F�b�x����<��k��/���~��-CY��B�'1`���xya�����i�	֮E��Y�&
�q-��҂4���tK���	�$�Ǣ���<cZ��O�_/��,����/�b���TjQrb�(�/\��1�, zA<�a�>�i�
�u<�`!�?�2@����:l��f�c���EG��WM�F�`?������"�t���Wd��a�~^s��z���~���p����]<���s��d	x��65A C��x�C��-�P�d6�y�D !3=��e�W�=�͟Y��9���>J���*..�V���X��Ptw4�W ֺ6jA�e�!�BGt��,�6�bHN��R�n&٦t�c�n�l��V
����FPx}�{���7���9�):X��W[�����Q0�����,���xk~{�O�)i�.;�B�$��wt���t�9I�bfe���i@Y���
|��ˆ��[������>�3��<@�k�Ya'Ƌ��)e�m �o{��p32�D!$�

/`$����@zm4t�&]]�,�� p����@�+�AMc;LJw�/�*�-Ǥ�h��oG�{��� ���|\`)���Wtb�f"��a\M���a��,���o$������c i� sq���q��� �]��O72��7�S���1�Qo��̇�zq!����@���֢.�w���J����nr�6rz����� X|�H�~Ɇxΐ,��"��O1X�rk-�L_<��e���1��5�&I��gھ]{�������"��Kܑ,����P"ƀ.�cT�cB�b~>qND�� P"щePD�T��)��/��N����a
œob*��DMF�Kҙ�N���B�$�a���=���/un��#Gد���z�Eӿ���DN�Y�阓da�q��X�!�||�=r��VFX��υ���=縉�{�*��ʧ�{�ǉ����l���a˺��x]Ȼ͸ҽ)�z7�L�Fx��<N<�Q�)�E\g/*I.s�D @����*E$ �l�*@  Y@��R� ���
]KQ� �Ҳ�{�Z�+(���X���q��M������`�v]�\1��#4�V$�Ѓh	G����bK�b쥤e� ˊ�#1��U�)�YFM*ȭ�H��V1�lH���s�h�\���0�lm��щ��`�;:S�]kyq)��Vm��+E�VJ��`�L	I�i���A�3�@���4)e	ZL���k� G�1����l��s��k�T��׉.j�.�a�ΛRL��;���X0QD�r��,V*h��+�y���D���l��PE fy7w$� �P*�x�v���Zg%V��:�asv9YMkv�.����B9l��Uzit��K��1�^q��Z�ʊe(���#�h����{���2��ؼíW)�X:l�7��Q-z�� Z���?!-����,4U��p3,U��V���\.��,�����m��i��"B9���q>�a��P�ʷ�"�aƼBC����e���0�7��=��7)�Etp�"��fmYt���茜6�����״�i0Us���SQ� �$B��@a� �Yc���8ʇ+ �S�3�"0Q�����Yhy�wb�c�L�k;����}����#-�&��ȗx4 ��R[�o=ˑ�1o1�!1�Z�T��1��a��zyNa�^ �O#�{3�B_�X��~�F�װn�nְo���~-�vD�UUP�ܗxN]D	BP!�"�K#���g� |�������(�y-��K> �-�¾�6ܚHbך7�@�K0�~{ ���w�.��}ޞ]߼�����>����]�)����b��������u+��1t��-�Z-��[��&��7$ �ҽlZM�k��[�Θm��7p�X*a+*�v�����C-dI��]n0Si�Y3�%�l�+_�	�P�/#��~�aШ�oq7�9kd�,���}M�̈1�� �"�Yd��}�s�{�>���Xڂ	Y��L��+��,ow��ֺ/��w�G@-�o3̀�A�����e��Ξ���3x�n^���&*"/k͌��\�����CrZi����/-���Nnz�s��9��h2z���ܓ�4�@�2��nW���|�O�g�&;����9��6��c���;����uܥ�voQ0����%X�\;�ލ����V�(��}��ǁ��y�a�����M�z�s�2J]���H.؀�3]yj	�ߗ�=do��_[SF�["n���L=1���om�;4�Kz�T�����o��D�DI���o�fo;�g_z�>u|9��=��]���s~�
���X�������p�hd���r�Y�g3Au�c�[ �����śYykv�iy�\71�ʪ�*�E���s��O��cx�����l�Ć�ܫ�J�5����x�󰰋yXpc6�}�j�h������lw��X�#����P@���]�e.�7���������9��7�� ¾��=�m�y���ZBv�m��a�`����r��5�2�&Fʙ.�K�t"LCH�&&GWx Nz�yv>���Y��ܫ���}�}Q��"Q�]�g�fx�O���6�-W�;����������=�vUҦ��bը���{/d1"ɴ}�1W��}���y�Bly枒)a��
=R���"}���1�V�$�=�Y�QH��1N*��7')ay�@�������򸧹�����EV�g�T{")��i�F�,�V�OeN<�t�$����+�PBe��>Н��$�^�K�ȋ�'��#����UB����

J�0�4�LE��1$�LI0LD�P̰@L2C,�X�,H�,�2R�$�ADɌ8b`�%�&!��q�	�2D�II2�11�.&d�h'�-P�!I@��� �'}6��<8iq�w
m�@��P<.|�o��P��*fa�-��Hc&ena�oޫ�|���O�<�W/`6�@ ��w���o4e�OZ~Ua���\��A��w^̲.NlJ<�������� ������c�L�|k�����Fm�	'�m��z���e-� B�40�H�����=�6��{qM$7M���=�� ��1�>���f�j���f�6no2g7~�Ͼ�����~�z�r��v5�"1X��Tai[R`�ژ�-�t؁&M��va��4f��"+���$�d�]�wnbTbR��I4���oϾ}��v@bI<��Xkcm��բug)ɰ�4{o��sP4y���,0�Lf����|�.�z�.�jR�1�n�X���F��y����Ȓ�NEՇbu����ڬ�p��j �=|�� ����=�X�o��:����V�]�y^w�VO�.J��s�E�K��D<;'xM�a��
�Ky�0�6� ��0��۲Q�٭y���㻾̊����_���Xx��;���]n5����nl̉��BF!��"�`�J*!���f�Cus�nkHe@z 73��tl�f� 7����Æ�������vR��ݎ��*���f�NH�7A����a8q���
��i_k�'>ϯw�󺮼�k.�x��+��7������Lݮ_����;�u�����^�K��1	�d]h"���ܜC.d�)QBf|�We�_o��©
 �"Դq�f]�8IU-yjGZ�$ƌH	t��֎��)c!4�'&��J&�5�n>�_<�X`=t�e��{�m����=����|��}�g��r �����C��Z������
d���nkm-o���[ g��#�"3A�Tn���'��ԓ�� �zktQH��W"��xt"M�6w��ꗎ͆徸��Dn���X�9���zx�]p�`	�d�p�p T���G �U��a��yO�zaZ=
�u��p�� �p�i�"-�=���Ⱥ�g:���xG��y6[��7W8��|���sk��LE�A�̡�ݸ�+(-�3dE;��Y�����=}�az���I�O��TՃvߞ�l^���� ���"�+\�'{7~�:��ӑn�3O��q���fZC��]��w/�ID?-�5�l��k���y����#Q�o����p³Hb4���.�-�P����#�{0h�C���i#Ԙ\5���
�����O�0  !�L�'� G�8��@tC�&:��O�Mz�G���>���	����N<�<A�
�;�w��7v~<�G���M���� L.m
�nm`q��t4�"4�+B&L�,�&8hk�Ĉ)��v��5��ɦQC:���!�P@ඕC$R@H�!C��0H�&e2�$@ü͹&��AH�^&	؅3H"s8�U1�q��
a ��k��P��E���Q�4�I@$ q !�l"��2"k� #�DHD����43ĠP�T
i:J�1N�����e�Vl��,#Ì������8
�.�q�p��C ��Ҫ���D���G̈�$H�)H��@�����SB�G�VNu�'C-�o��<��8����`pp��}�����	�j��1��^O�W��͌�'7'�#B7��B�7C�.�r�1hq3���;a���H���O�g�Ɓ<���eLs���˓WZ���DUq�F���{���C��?������&�㧫}:/%��o����@G˻����]ǁ��> Qr�����^M��*|T �w��"(��8���0����z��y�}��E�y�~�gq�l�x��uE�����@2p�s�G���'���#1�R�蘹����O�7��Aؠ��"�#7r-�f�����G��uN���I���(?g��M^����O�ICD�ǰʡ�'������c��͙L��M&���)���� ��]S}W.Wd�4OdG_���Ǉ]���1��L+�<�����s������R>��X���(j�@� �!z��8O����� z��?`H����L&2q�4ۦtE7*(T��0,� \��f`��U�1��PB�C%E��
�*���hF��(A��HX!�	s	�%�	eA
 �Aa� e!�)B�ZV��(A�T�@D�TA�@BYQ�` V	XahbX�a���fI8)��)0�ұ P!0�@4��EU(�
�b@Ċ8%D�n:��$қ�)��(i���F��+��#����@�	�����E��a��H�����8�#� ��T�@�{�������vv��e`xw��G��/q�9.����(���K�y��s�x;=JBzʘ(h:����>��<�䟩�@���BIC���S��5����E���t[��z��/�`� ��~��1u�� �|+��+��J�(i(i(i)(i)�JJJJJI�JJJZJJZH��JJJJJJ))(hhh
J)e���)ii(i)(��(i&��������)e�����������$�����))(ihi)(i))����d�������	)(i(i)I���b��i)i)$i)(��"I��������!$�i(i)(i(h���ZH i)(i$��JJ���(fH��H�!��i)(i)(����(`�����b�����$���bJ(������i&JJJ
JI������))(�������������������������)(hi(hJ))(i(i(hi)&))(i(
�����JJ��!�(i))���
JJH����JR$i"$��))&"&H��������$��I
JJJ$�(��ihi)hi(i))�)ii(i)(ii""JJZJ�	(`��������������d���������������)i(ii(�������hbJR���$��)(i)`�(bJ���)(i)(&H��������$���a�������h�)(i(fZ�$��$���ii"���ZR�$����������i"JJZJJ&R�JR��hhi(��(i"�!�))��������"H�b�d����bZJ))(hhi(`����I�!�(
JJJJJ���������������������%�����(���i(i(hfJ"JJ��$��))""H�����!��������%���(h����hbJJX��JZ�������Y�������$����(i"�����I�������%��$���i)hi(h��(i(hhb��JF$�i(bJ))"��%)(i(a�����(hhfJ"(i"JZZJH���������(hhh))(bJ�*�&�b�(�(��� �!�)�bj��bh����()� ����)��P�������7ҞR:	��IuA��h���� �� ~�9�쟚�S�1���qW�~��8���8���9�tɹ�n���w�:v�?j|��W��䯑����y��q�]����)�	��_G�M���}i���ɪi�ԯ4;�c��c*���#����UP:�ҦҞ��%��paI�R>���M����N���]v|̩���˕������=�`z���h�������Y#��@��q>| l.1�"���� �}�0�PQ�ژG�c�Ǩ^�����44uO�'y� uل6��WW�`�B��4�2����ɃA>��'z꧑�TP�e�u�w8@T����*5��MU#t#�������StS{丨�/VN�h{�bF=������;�N�� a;�,�q *qN���+.4�(vq��N��#�p�w��d|"����X�$�: b5EU@�&\�¸1����n0Bz���A��P���� ��!�������M����G�T~���ہ������f4���+��6���N� 1��@_Bn;��~�Tԙ=P�`�zS�'�q�����o�����%�'a� u/D�8G�G��tʨc����*(o�7���?���x���'��U���=�{��~
(�!bX�=��v���{�E0�����v�������X�w�:�0��li��w�hn{�ގ�|�r������Nr/��^���8k�D`�(��x��H�d�ӹM�v^�M��|E�	������]4�8��@�	0"���p �팇�p�Ln�CT�h�jib���{��G���=OctT�c��;��0hmd=BzD�M9��
����o��x?c�~ �v���&�� ��:ta4Gq!7G��;��φNGRs]���W����XAMP�L��8:����O�OBn/�t8�����D��6��4uN����B�/���?�`yzO2U�UA�Ѩ` ���MT���@}a�"�	�L��u�]��j{ߐ�9� #�/�	�/k��	��u,A��_jꡞ�nq���+��xr���۾��t�����!�!��kN�=�d�7tD;���ǇQ/��!�cP7��(�����)��3�