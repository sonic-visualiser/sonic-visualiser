BZh91AY&SY��j�	�߀ryg����������`�~         ��z       �  ��B�P� �
UD���(
��Tn�ڳ[^����;�K��3�h���q@��ܹB�>]��q@(Q�޼B�<  �EE�\P
uw\Pus��@oG����QE�\��������T����=|_g݊>٫����ֺ<�N �Z�{���Wu�ƅ c���;��un���)���(�E<�8������CR������47N)Ѣ�β�{�}L�.Q��j���P|>J ��
H            րA  i�)R��Sbh��h�0&i��h?U"2�OR6� &�&F&F���F�eJҩ��hɠ 2i��  a��QA)F!�A�@22��0ba
�&�1��2F4�LSS4&�zOOG�A&�ڢ	*y�SFM@�4� :ǳ�{�Ϝ�|<sx" �����T�?�B�D� �AK���jDG���`(���a_������{o����4��������������]��2����:.������s��m�\���EBv�!���Ʉ8�AU@�2���UG�ĩ�Lb������я>�dA}�q��׹4E4B4��� v6z2���j����s�Gd)�<s��I�0�_W:2)fu�zR) ��B�� }�7���|�Zcs����x��?T�L���dя��{>��޽�N���|�o����nB��V

����ݡ�B��P���V

AA`��PP�!�T���0PX("�ACAA`�VۡnaP���m����[���*������A`��nЬ*

�p+
����
�AAT
���m���j
�aP�,*�^v�+
� ��PP� ��PXb��з!P�*���AH�P�1�-�B�PX%�B�XT*q
 �P�
Î!K��
����
��¡PU���[m��(V
�B�V��AA`��\AA`��s�X(T8�0�V�q��k�9�m
¡XT*�B��eB�m�wv¡XT-�o!P�cP�x�B��T+
���V�hT+
�anA�
��9�T�m�
���
�aKm�Xc�T+
�A�*5
��C��[m��B��
P�+���t�H=b��\�A`���PK�ơymݡKmݰ�V
�m�
�<AAaP�
 �����B��V��[��۷wwwwwwwh[x��ID*�B��Pn~s:t�L:C�+
\
�qB�*�B������B��[��7����j0���
�¡XcP�V	������!P���XV�V�T3-���uCXj�B�XT)p+�(V���(,*o8���A`��s�
���*�B�PP�*C�B���
\m�B��TB���#
����a�[��ۻB��V


�A��� �P�*¡�����[�B�*�i-����:�!����c�T+
�aD-��*�o�PXT(�V
\�1aP�+
\
�B�ơP�4B��V�p-�Ơ�XT4IP��P�6����p+�g���*v�hk���B��T+���*�B�*
0�T*����Vp+B�U
�anB�P�Q%B�TB�XT+
�B�nB�
VaP�*���r�+�aP�VaP���-��*rC[��X,*Kr
�B��C�*��V
�p8�0�V
�aP�j
�P�*	p+
�Z�B��VB�VB�_�0:C���wl*"���B�-B��!D+m��*���m�wh[�F
��Q�B�׍�CX([����V
s�q���aK��,-��7w��A`��)1�2T�"�Aa�.K�/�p   _*r�d*��e��~��y�>��w�s����'�׮��'̷���d��_WfI����0w��?�y:,���1{m��m�{`˫�����4�>�XCɛ��	��pY!�ْL����ҧ�̘58���EZ�'.^��zw����T-B��17YN1�T4���u�Q>�>��б0�DĘ����Nl\��)���8�&qDý���\��CJFA����B�97&�.lڜjw>�_�izo}B{�~S����>P�yQac��S1"d�eϦ�y���*#��\FK��3qhU	����$[aqSYt
&��ӂQp�˔*�2&=�J�"��r"�a�[ϕ<z(��N�$�쌑5��x9ʺ�f��<����ɹ�Th:��MR(�J�T̕�JURǊK䉼�J4&�sK.'�/nב�l��T�"�T�����D�����?���ȧr*���1��S�OT,KʇY��2�2�2�&'!苌�����`]E�Ooof�h��w�9eԌ"bd=�9V�B��7W�f�v�4�HMAs54�!N1P|���L�8��w7��Q*Az/)K�ɂ�E�6UMӨ���pM3�����4��+ǧu�P���sj�y��*.�:���8��ޖ@�#&ng�/Yh6����E��O0n�"�32b��|�b�9)����1Ɣ��ӽڋ˫Į�:QO�C٩�2bތK�H�Y �Zz@�5Ug )D+�Pb�AX��]ԨBީ��
�Q�E��=<fVT]Mh��T\㊣�H��s �\�Rf$@�z/�Eǒ��D=�J���U�osr�C������Fd��9t�G+�5��/�'�1QR4&q\��-D=��H`�U�UH��,�B`T��r2���Q)'x�²�"�2�Q���^3"$ԐA��x��iUX��ʚ�F��
 �,��13=͊e�Sp�c.i�Z�y�$�"�J_O�y-
T��]�|�@�M�LZ��̼C�ʅU`���$�J)��U��sX�d("P�P�8�9�T�PN�SR(:U&Dc�K�Q�e&s��j���e�T�."f��($�&*rU�䨌�r-Ռ�����FRʏ�p�c���*2� f�oe��u��0ȻʁUe�%�}*�����c$��^�7�qy�.�ګ��/��AJ^U��6K��x�9w$�Eڻ�e�J2_1��ENMK���7j�Nr�$C��]��^�.U����U*�q��"D�
���.�ȥ�T�QC&r��/�q7�`/qfz���A	��B"]�BI�����wn�r��l�v.^b��S¢rc#*��M
7j��f����L]��&��B0UʡR�xus�{�r�T��4�POO*���Ǻ1a��q�^y�������ϭe̻�s"c#���2�Y%����ț��Y�X,�cҩ
/0�e
�)#D���ND����pf��T��y�˙Ȝ̉L󂲢`L�Yw'2��d���8�b�ȫY��
�Sq��K�HS���T��e�HU��7�1.k �̽�*mI��������E>C��(SHS�s)��^]R/Y"�e�3�lA�Hc�[��N�t����U��B��E`���T��MԘR�kQ1w	��<da�&��J�U~{�B�3��^����_|���||��i?$��waU�U # @�q�tI�-M	0�PK�H  �`)[�� ��4 H��
B�� Pݩ��  j�Q �-
P�+*b@�ՐU Av��IH  
%m��� ��C%n䩷"�X� ���Z! @"��� �]� 2ɠX��,h@"�P.�d RHƂ۔����(�p5pP3
�@@L��M9!�fAAdlX�@���4H A	��]���L��i@@p@p�R"
B��Eʸ�v/qX�B��U����&��������5��m��3��ؾ�^Sؘ�==7��@�:7,�1�>^;�x�<��������.8N���,�;�����Ӯ1mw]��]�����˞�sL��3$I?ݱ���0P�L G��%R�n�0��[��JO��X���W���5�q[vàa�@�	b�!e���D[*\^�k���xF�V�b۰�m"!6x�
�r�a�L$#(m��Le��4.�F�%δII�f��si���v�8��,�}S��M��i�LC�Vhʥ�y��-B�Yԥ�ւm��@c5�?���]ې�T+bY]4�� ����nH��ؔ��j�k*���B��#rS5���MQ�ĉPv��$�I�R�357$6���e�7.F�!3�KVd��l%����Q���g�)�]+f��u��&6eUn��Jli����л�CgD�6�4�)6.�Eì
�0-Ʌm5�����.̴Dִ�E�4WY�Zmh��]x|��bR��]��D"ͬR�5
�.İP�j1����JsR�N�A��5�-����y�6�йa6���m�±0Vk��jB�Nɦ)eu A��=Nak�Ue����:5���{d�,�Rڌau��݅,v�(l�X�f�]-��2��������\ۉu�qA��12Q��hXfm��\��]l4Gf�lQ%"z��z<Y��X���]3B�VhZR�WCkB�B�Z����-!,c�E�n��ō�Jn)�ݺe-U�k`�%O;ǭl�GA�c��e��fW&6`�"�KpLgh��u�S.m�[��!��ek�35��t,)��nm�·i��`�5"�^�"�a�lmN�a����h�
Ya[Lٟ�|�W�B]F7-�hGIf�Mche����*ڐ���[�j�mZklcBxl+X�����7-e�%�Vͫ�tܥ����Gi�5�d���`�[�NZ�)�:Pd��^l��]nd��S �; gf��P�1�of�Z��T�F�v�5d.�4�J�e�@�%����l�\J㍔���[�m�l�� 1�]��\\�fm�V���4x��!�&�!�e�vMY�-�r�-�,�d���4�\�����.f�V!�!Tn��)��H%@�\J�#j��k�@���f�z�e��m6t�+,js����;J6�&,&�lL�s.pb�w3m�f�$�,v �,u
��kI�O.�zuv�d1�o.�6�3���� �{����7��u�DC~��<Kz���=x�U ��?�� �:7�Ń�G���FnG{�Nw����yCȎ�|�������~r�\��8��{�/tW�I��ݾk8��9�^08s	��-re̊5���ֺ�s���B1��F�<��;$�<�6�I�Y�=ou^����e���I���Ou/o�C��	�G�~>��u��)m��OH�+ �����=e�2e��+�b�I��+{�}y	�o|Vy�q�����ec��j=aY	��p�@�4��Z!�첒%�{w����}���>�C��=iy�X�R�#Y@�x_���������O�����{n�֐<�N�Zߓy��s���{�f�0�jn*���L6�8��3�^U���X���ޣoϏX����eP0��'�@���JL�eͽ��|�S��Α����ҴgS�h.� D�(�T��y��&�ZJɧ3����H�-����C�z�`��ȱx�{x�-�e��B�
u
��a	�����d2�L�5�33>恵�]�ʯL������R�&e��T�R��^�Ni�(��~w����ǧn��/&���צ�p�<L���1�%�8�!���ªE[ς2�=�L�&$㬁X�<gt�`��d��A�hpJ� ;�Q��>�+(��5��v�,��hwU�s̅�b��̓�d����|d�$ C�˯DT��t�=�u18���:�CǛ<||
}m|���'�_��l�e�z|Sߠ}�;�:������Ut�,�#�?����<�&׎}w�xm�=&	D�YU�(�1�Ȱ�bҒ�4k
P���R�$�S�!}m#(��>}V|��@� F��'˭f���~wש�mv��C��:,�������r��O�[5C�l�yD�P!#Fji���(l�=�0ЕӁ5h�Ż��w���v��LB �{o�k�z|��%̽�=�ߐ�;˴�r 

���F(p �X���=�Ik$��N�yg�F�����:56��P̴�cd :d�9���A�f@����� X\�;�:`gO<d��$��fzt����:S�#���Y%$���'���>��$�gzw}җ3��G3=&�q��C�s��!�gL���t��2EK��J��3�Yu�C�ght��=O�e$�Jt��Z�=���7�!�p:�9�:���>�� ��	$�@H�@5]]�s�p�ք� ��T����?��!TP$�� ˢh5d�	!��%h�!�AX`�#vn��@ 5h�dPM�Tj��u2]m�.�i����ɶ�;�����c	}h�UR)B�5e@X� �K�&�P#$�����MUZ ٳe�@]���]Ȓ"(��q:�Ȇ����B�!|7�:��s�ny̳lE5��p��k6W(\f�(#\<'tgx�@B�pLl�֒�o4I�D&Ö��E����6���,
�)�\8�S�[Y��͠4e�0���-�B�`�ی��t���SLBƚ5"f�0��AAΒ��SUB$7%�86�4�e@��G� l<fɛk�h�(U�
�2X �-��f�{�jR�ؓM��-�ȱ�`ib�,��k�bQ�wy#$7=M��58�Hk
�)��ҍ�"R�a\IN$̗(`��k��E9#��ś'?�NR���{~U`�PB�f�33̬��%�l�a�B��y�9f�9��i��]��wlp�ܶ��h4��)�FbҰ�VE9���m�����3j$��N$�6PK+X�����?,7���q�����v�ث3�擌I�i�oW�65�����8--�ٷ�b�2�*I'��a��0� 3:O��ty��Ś9=F�\A�L'>*=D�h�r��>�7���:��^���kmm;e��'��[�o�sw���ɔv(�5�y�v__p56��>�h S���׷�cA�O�/S�2A.."���yn��o3�����m�Nϛ� >�(0���;�5\��Q��	nȜ�ް+�Զ��W�����憠<Ո��Z�m{b�$(ާ"3�F]�z�Qi�z����Xm��C`gSaJ�A.�x�ñxx;l�1wiz��@���w^�=4����1@z���^T�wכ*u�M������p�B���������\�<�!Q�Q�$,U��wו����������ڍSl[��]ˁ�3�l��O7P|B���V#&Z[e���V� NebǊ�*"�N��B(������A��۸V��}���M�b���f��٧t�m�� T��<�p���@1*"!@w��Z��]���T��#��rv��<��Q����4	����"�٨��l���!�ݿ9 ����}��l��i��b�2��	言�!BO���D@�z٦�P�mL<���C�%{azZ�Q���K��z�e�iuE��Z#&#Xy����ۥ�kא�6�2��vGV܌�2#��/!��o�{���Ml;z�G����_�Lަ-��p)����m/5�/kь���@�D����Y�ճP��<ʅ]�"� ��rR��Z#��n�z;m[Noz���zZ�
�A,k^U0������jw'+�|��ky,�@Չ0��D@�J�סq$� ���I�S����r�O��� W$jIh!vt�u��`��Q�bX�R��z�g���(Da��B�ٵ�ɂE6˶)rN�#&�ݳ'#��	�� �X�;����x7��,��i�1�ik�ئm�	���oKy������j=a�ג���7g{�9�2��-.M�p���尶C���O��=#�T1R�]O���l�����]TTW���f�f$�`�� �JXkU[����-���P����L%��b��m�h�,��e�a�jk��$�L�9�M��s� kۍ��vd��ہ� g�bA 7�f98��d�s�Җtk<��p���<��l��K���zP6�EJV�+��&<��R�.��=>p��S���/���SG&n��� �3燤��#��QJ������F`@�_�#0T<�����X��%
�[o/��FX>�"o�����11���1��v���Us���z�Hw8"|�b(�!�}8s��L�y��ܝ���Y��g�{z��� |0��'q'�d<翮@E���,�ɼF�u�D���+���Mu.Mݖ�߳�'��8�;�7����k�r'�<���	��M���m��6ŵ���U�� U~�zyÞ�߂�61$X���y��n>A�e2&@s�<:x�"	pK�0� W(��c�*�~�0�[J¬�l3����BC� m�Y�[87\�T� ٝ,ҵ��Z[�;Ⱦ����ެ!	c@1��ܣz�h.�tQ���u9��d@�F)JMZ�/Y����nk+���5�F4ѥ-]�	Hʳ�E�A��HRe\L_ս�@�kf�����G��A҈xxv� � �h
���rA��E��v��8���ڰ���=�fX�����E���:���2�y~_�z|�cϒ^��vMh����p��3��N�M؄6�T<�rD�˖�K��-+%�c5 pF�&�'��
tɶ q�#ѯ�l@i�n��mm����ۈ�*㹠 �fC�0�üAxFC�&	)�Sx�c����0=�� i�e᧲�@�)��:��D��~~��{����jc��&za�8��|l�y)�>b ��c�]/�~K���0�U��Gz���,�=P��v�ɨ���揭��q�d����v޾p( ���Qf�&
�q6ܤ���q �R����dL	޳^$�` �8��n�膖�5�H�Mg��Oh����tn�,bg9��3S��������;�}2Ȇ��2�?|�l2��evB�-&�:E��;z�M�* �Xͭ+9K�!�\d�>�v~""& �ALλ��S��ŷ�|��w̿qϜu�J��}���q��$P`�91r8�^d�"��j�Z�45e��%�"�r�sNGW�e�Gq]7Mu�Q��ͬ�2	v�O�{�|����@	!�cK�Kv0Tt���xi���:Z�xc�u���Hk�,�hlS����#�`���r�jG?A�T�I��;���O��3�\�õir4����#m��Ha�q�<@�G=nr���yf�a��gl��xD[ ���`��`�L�Xm2����c�N�g�#xG�%���;]�j���ͫ�za�I��\n�<'���1ӆ=ĉ�{�%�i��L�އ/R�;	���=�>cT���}���C�~�>ɩ��&�mn��@i�=�p&i-,��u#���ʍ���d;��"�)�����#��Yn"�:ռ����b��k鸛� ��c���Yzk6M�ˋ�:	����G���[�G?��仯lAJR+"DT�YU<* �4���?�}쇞�
��h`�������p8Zx�]�6�$��l�����H��C@omgBTĦa�X�(DX�Ձ Q DE��1�J�K�
 �1B��=�~�L����tP��/_�2p\,{�/19�"�Lх��g�.���k�_���c�C�LUD !@�	��"j&�2,{�TV�=�AJ�z^��/V�f�[�z#�aZ��A�W�6�;��|Ǖ읬���x�T���|0�=OY驐��J�>����'�u�������u��ٿ>���� ���  ��/M"�!H@ \ AB"a��&�a���@գv{S�ɲ�˹�]aR�ê�b�*<&��ks-T��c��[�Q�	`]���1i�M���K7{Յ٣.����g&F	�˰:ʖ)i���b�%k�h����ؚ�X�IJΘ))�DԴ�C6b�6�6I�͍�l�SDU�(預�K����5�)Z�&H+5jRb����R8�GM��-m�5bl`WKeW\�T��,qkJ�f]0��l�sGQu�v[ͥ��X1	s���7��vO��⩗�S�$۪���Ͻ}5D �6-y~��毕�B� Eb�Q��u3��ҁ�H�bb��������8���$;Y�rX��F2[���<�4;�׍�X<���-îK�g��R\N�ﴦ��������k�io�5�H���-9����t�6i��Au	aly�0=Ʉ�C��y��-2p����?�I'd�Nu��j7m�#o-U޼c,���0+.<��yZ#O����G,��uE�]�O�N��m����[L���Yc[F�=k�gL
M���;�͜,����0�~��LI��"<C�(�D"Ix��"�H��a���r;4cla�su�:"t�A������� Y��і�Lk,�st��q�m7qc*���$�at�[��c�,���;l�v��.h� t�(:CI6�[�:��M�\�i2WyĆ�$�Ũ�Q�oC�6��
c���3������c�<L��ǟhӀ�\\�����}���
��l-6������t�H}�Ӿ���<�4�2��� qXXX��׵�'�D0p�o{�KqƶZ�WʿgU^��"����Bp! >LC/j1?y�P��h?���KC�Z�*!=$3��?LÍ����1V�gU�[aD�[Sc9�D�Ƈ�> �x�@ Mz����l��V�r��	:Q؇w���(�3YY��%��:ű�5t�IY��d	`�Jy����� l�2���xr�Hu�d����Ϛz������\2�DOC��ۊػo_8��'�Y��<]H�ɑ������8�*����ky�:�L-�p%�e@�4�K��cٞ Q�DC�l�A�D���)�)�%	��3H�X��adl�Oc��`A���d �Go=��2Ǥ�y,ʰ[��:�,?�5�`�F)�8t�G���di��mc@�;nx<�̈N�;e���U!ۼ����}���xi���8Z�����1-�U���gX�S������9e�g���n^�B`@�ѧ�iӭx�fz;����cr.��a�z��6xh1d�v��tD�4wA0Uk�a��j��A���O fS>���5=��}�����$���JB!�"fF�GX�	
��x����/�/�AQ �Y$o�κ�[�_f3S2b�������1u�]l��Y���Em�qaF�˰�,�>;��eb�k��11흣UI=�����/�����+��;�-f�r�3�Z�6�Y,��唦�U4����<��[�h^��9���,����dhic�̓a����t�(�8�n��������	&�*��Pc��^������
m�ݾ���,�;��\c��K^�gX�>�~q$�-�� K��1�fd@I,�(gTeSה4痟/�S�{���&�4�����Ǒ�KJ ��	��K�a]T艩�u�'��E��^��7Յ~��W�����_����V����{�s�n�����%�����B�Gk�~>�:���!D�p��y����y��S�c���k�8|�P�R��2�
8���H��dy>z�գ��[댵�K����F�'�e	ʿW�(��0�U�v�N����T�����	��	8��
�EEUR̅P��E!��ERTDA �"м�i& 8�a;��:]�~w���3�5�a��,<��?�N��E%+{�1S2"+�
��̊����쟎<�'�� (�i �=��@���XTI�?d� Sb�Ý�#���	�55�9�a9�Y�ݬ':Lb[F\<��	�07{���/ٴ��cqC-h�+�)DD=(�Æ��27�VŴ@�F�\	n4oT¸��ljcXb�Or�Q-�`���a�6_�DDD b2�XQ��sۗqs�/�%On��M���}޲|�@5p �gؽ��]rUh4�Du,Y�&�,2�=GR�V��uռ9���%F-�+�*�e���A�Y/[?E�~���m��i�ei�锷�t��gM� Xo!vC����[LZ�F�C��8�����	�z
fa�E�N���H
"
��i�Zϴ�%w�Kq��$�D!I�
�x�dD8M)�=x�w%�ǌ���0Kw!GK= �{���1l�Z	"�O�y������ĊD0Q+��9]���9�ɽް���4�a�:�����h��a	�$ĬNoUM ��&��=�g����Zǁh ���߄��e���0ۼb����de�D�v�a�A����Q� [�OO $��d�tقӧ��y���0��lw�z���f!�(���0�ȱ���f��s�h˧ב�l��le��>�Vq╢�c�ۓ./+W s;�
,;����Oc(,��N�,us�inc@F�����xj����}ݓ,�cLMdL7���DDZ�P"+|�<�2V^]f�:���Y9}�\���>ۮʃ� V,":����-]Q�vu�m֬���F+	U�mR��m��塥d��;�@�kjY�١vm�+t��;�}�Ӥv�ڞc�)��Z4����Z�d	�7��ƃ�00"C�iw	n4v�|�������(�����Bx�55�2���L"[K���PDv`��;M>q��ct���r4��nelCk��ߝ��Ҡ� Y��W�:[�S'�ܗ^�ϋ��(df�vm��C� 'xv�bH�۬��%� vHZ�&W?8y��LP�E�a\��9�����&3��z��Z�!Dx�E���x-<�`�ٟCw<BJ�Dw�͎Ц��Ձ�|��2I߈~O�� ,�-o�M�2��:	"`&Ѧ�xѲ�p��{)K K ��(��~�O�Y�o!�l��f�-	1x�q�l�yg�:y�����{����S�	�y�h�p~d�cþ�@��y@�p�~?s�Ķ�GX)��[�?!$��-'L�!�;���t�T�4���46>���������Th�U)��s��-h�_���8H �?���s" MU�"�ݾs��99�(�! Q�_|�9� ��\˪�?��g�×������A�3��ׁ�Q��%�<D]/z�քԺ�FBLaqD�z�$�bL�q	���'�bk�ѻ�9�>�z�SJ�=Va�2*�z�`�x�u颭c��<�N�x������M�r-�� z=wJ�n�-Pzx|�|�ȃ������Da����uV�����-/OWtw}[�;���Ub�E"R��P���f[*aJj�B�EM]�AiKĹ#J�K��FP@j��DLFB�Ό�g��K���ղ��E"�6f���5L�ms.�[��0����n�n.�mE�Zg#���nH4�r���F캮1�ki����vF�!�LM,e�ٔ��GW]�M×�`���.�27\�۵q Rƕ�D�+����7+*kF�^h��i�v��5�.������@hV��[e�B���r���e��V��T�ن��)W*�p2�L�b�V���:U+����xoY����`v�(�)2q4D���
Zi��(��D!
R�j�$hJ)(1	��"He�PU˻�r��o._�w��H5d����Qr�m�B-��X⼫�_�3��vvX�h��"�0eJ��%�5! ^6�@G�Ts,��
�7L�f
I�s��N-l���p*j�b" ~r`�&���Di��?:x�_|�4���i�6�D�=
a�`��(�x>�C���i�Z����x,���pX$���{��>�~@;$�\l5T�,�;��@38�/�+�L��z�����'�D6{�S��A�|*�o��Sfkٟ�8�Y6�Q�1� ݹ��[�q�.Yhq�5��A���'���]��0Y�l�2��z�e�kl$�u�%�Y��!O*�O(���T���P��V�lm1�+ =���0rt�5� 6��\�-��r��ɾ��񲪎f0Q��*DDCC�8����lΙKy�Kd�����|M,�	��"0 �l�~��)���=���xlqƍpi��okY��l��jsʿ��>����^��d��2�njQ�U��);϶v�	���Z�Ϩ�%���@[ϗ.Xq�`-d&�_	�gkjR	2��z	��倀
��O/何�����0�"��"!'�W�t�_��BO�2 �B&"ah����ޭ���e������G.G K�Y��%/���S�у "!�!�f�39�eꪚ$�]�����s��##���'��X�pL�@�Ot�������{��c����~���@<���~ˉo��Zŭ�`w>c3.��!����TBpΞ�F�w��䫞w�����$��T�,8��<ab�l8��J� x�~y�&��`b�or�ܕ��_WS���٨ʙu0�kL�����='~��y|��O'�R��a-�pL[K5�;�=��Sp�PpXӄ,�������E0;�y��-�V����6�K�\9��>��f@���݂032!�C�>�W�7w�!�.��60�<��t喥��!�`$��3�v�2��j���5�nZ��;
�#OY#�-8�V��&׏`L��B}y�<��.���Q��Q�%���K��-UU�"��d����W��C#�i��6�$��i�r�����玖�4�`v��vi��Im6y��� � @+vlј�I�۹�}�3��;���Ϳ~�\���U���mh"�+��[4��FX�֚Ԯ���6b1c-��k6���Yo&�?���P���>�-�.�N��>����� ���f� ��D�!�i�|q-Ŭ���۽n�6��@�Ei ��,�r֖�7pƃ�K3"I&w�E9*""
�10g�Z@��4@��ˁ<hn������2�]�HrUx�ˇ��K��`<��M�8�m0��WSȐ<n�^b1^� *fb!�<C��;��I҇N!<@�!��~�ޢXa�l��[~ ��������y�7��"9M<Y��g���yo�+�Ij��*���`�X*��p����j|>F�<c�b������4�3��Q.^1I��o����yS���<�(�m�FFO�ytb6��t���
��"ț���MF(�371�\y��]]�V�_�����$�E
q�(܀�c�{·Q)��2�Y�U!T�E�CKCUEPPDRҔ�TE1RDR�$CHR�R)P�LHU1%@APR��LSSMIH��:Ț�	�*��eV�lo��<�r�	tO����4�n���@����*�V!9n�OR@x�&t;	۔�!�"����O-c�Q@{o�	k����$w�C1h�� DUz���ψn�ya[ӂ+SU�R����BN'*"�Axy�f�"�� ,���'Ձ������A�1�6a�+���8CI�v������i�-�h��ӽD� ��D�fy.�r�/$��>��'�'}F{����`�"("�H�3L!��\��F]�:ْ����H�S����F[l�h�vcE�UUp�K6�Q��O��<>ϣ�~�z}�*�O`Y�����눉�U��l>�Q"ǂ��]� @枞@O���z���.�"2@-�+2\Q�Ww�w���el@�&U�8��G����J'���ʽ�ZN���:��Ì�P ��s���P[��d��Î�Z���m�fdAHû�x1��I"���s(�G��z�a�Tt�`\{���1jcC������Ϲ�b&�T�{�=��ahpO%�'[U�b��r��X�Dy��^�p��"D�<:�t25��f�.�޺�o��$O�-�[�P|���	����x��gͦ��@"�����v��1��L� �V���yl��d;��"�N�.����.�[�� �=�=$���?�t�$i�	�E�� ��C���`��2x� ���U�'��&������}��V 3.�
#^�a��LM,��^�ZHo�x����"�x�ĵ�y��8֚��� ���(�s���&Q�H����Z���1mV2mTK�ZP-f��Jm �OBg �Z'����$Z��N���`8 i���˟p&R�3^ME��� H�s�q�@s:4�}���ʪ5n��7��Q;9'ư&;��[\��=��[o ���*�k��qŋ����	A��o�����:�Z���U7&d���6��[�'������'��O�F=�z4&+ve����En���+�%}��=i�>��i �n���je*�o8�nP�ΘY��V�t�������v�a����1o�X�+�<�b��-���M�~G��y��3k���
b)%�DC�U�T��)� ���q@P��d�Cp�޷�«��,�ɗ����˿d�0�J��0�AI�.�7�ˬ뜋ˈ2r0l1�.�`ȡ�L�l�y�C�ߟ�]��.�����P�f��a���  �-UŁ�>gTX>|��E��O	��2�9*e�.@��xoe�����h�[��b �+t�Q�t�@Y,kV ��2���5d����Y1.�cP���DDDDsY{w���d4u"b<MY�5�E�+�TO4���5jZ�]�x���:/"�xx�t��((���E2Bc��|%�0:0���_yˉ��}�'�'!��/O��D�w�J���D�z|O�%�Le*��D엊U�<�	b Ȍ�>y�!y]e�
U2x�#��^�>;5r�үU<�֓�f(�J�,U���WuW�u&\�Xش�� R�kZ��Ґ(�L�KF.d�v uaB�1a 2�@�C`n��:Nusy�mJ����2эe\A@R��KnԎ6��S�5#�.J�;/�ĖZ]�ٵ�(�,�.�W,n�Vѫ�
�`�ˮ��U�L֕�VT��ƹ�ԃ�ٱl\˪�cv��+5LF�ċq-p�
:�e�[r1ɛfnS:9�(f�Sf��a��I�%+��6.��ͅ�X;X�Z��vz�k�&���o(��EJ&[�f3em���lm��1������t�$P�c!:Lg��,7���wwwtA�a�b��\�^Kh�� �"$�2a����kosI����َ�0A��V��%C���)"�����J{�ӝ��a��7&3�N�.S�k�!������z���h:l����­.m� Sr6����ja$i�i�L�~yԻx��oG�^󳳱�.EX-��TĴ�¨<�N�����{�I4n��� �<�+IH�Nי�� ZHV��gͬL��U�vjŦE (�S��s�KQ��BL�""�`D�ww���Q
��#�l��|'X�������	�v���OA��j�,zh���-�0l���S�4Ź��'T���KHS6�� B���"��@�ٮ�;��O9�=r�yg߾؉oGŬ���o�)�������\��a�e�Vt�Ф���6/c�Y�a���mS���8�bv�4Z"!��G*:�AZ��a�9;��y�τo><��d$� 9@�y������`���@i`�M��2����k��Ϸ��g��A�A :q���,�`�r2���>C�4@Xڂ��ՠD�jٺ�slp���k�;l\��.ɂbdf��޶2���F;lrI��r,��*�2P�"�	*�9)��h Q	��jq�&� �j�M� �kx�6[M���� 1�)7�j�R4���gy@��C�
�a��hە;'��9$�K��^�:}�H�YծЫ�eה���0���d4q�\Kalf,-��WO)k:Z�ah	�%\��a,w��_c����{vQ+0�&¬eՈv�-ne�#m���oc.���j�����p�ݺ�ڷ4��v 0CL��]8�n]I�E�g����o'�Ͽg�Q�.�gU[�a��h�YR��5�;��m�3kK!����<��t�b�Z���ʀ!���'���&D`K�{�*e��ez�?[��Ҹ��ߞy�,�4�މ�q�� �v�^"�� kB���ik��ǣ��0��gŀ>X�m먖�(��F�o9�+�׵�|ڙ�M���f���L��n^��%�>���7��u>w~w���B���zۼ�V�ۘJp���ֺ6a�-(2�@�l фX��{iI�;�w��i���&�!2&G;Z�w=~R�|��������1�6�;mo;O�A��.s	v<��'L���	�6%7����c_9�^�#��\QR��8��>�<�v�n�y�q��;��׊��v�u<�q���@O���!�h���D����d_�8ǈP�������<����>��/>s@�aqJʲ�
�DC^"3	c�l�Z5oB���{ 9b��{yoZ��N��9��O�d��q�y��ȳo�Lߤ���UM���I�N�f��T�.�y��<���9r��3Bf����X�2_�*T�=���^d�+�3R�0�y�^���S>^��r�I�겠ʬ�&�dǵ��@;zV��U��e�=��M�gRWaLb�9o"�<\F�&�xzMOZ��U���s~q�#*���}�J<�*E�_�EM��
����:�M��[����G�Oq-�Q�1��hB+�5S5�-Q�V�f���Y������>�3� [m��i��F�-0����hMN���u��m��bJ���+�Sj�m{��	��X��� ���a�`�A\	;�o>Y۹�����'�;iσi �=�"ȂNy��7 u���-��O��]}����" ��ﵲ������󯗝��}f}�'��D*�[�m#�9�0:�&l-��T�u��u�9B1f�5Vv�[Kfl��;�\6(���n�e�g��N=�7��e��o�Xx˧2[Fj�y4��7�Qmc����9,��\I��8Nͬ�w��E�3"D����!��wPa Y�<E�9�2k>�q o]�q���+�W�*z�k0fb@�v.�K6�bi��l&�:���KIi������Y�u���~y�ޒ�k4�h["s�����`�{����j��Xx���`���-=(#H�<wD���Бo�O,z O� @[�1p��}��_W��V}�����1��Ъ5(�5ΔC���`Z��= �K�Οp4܅C��D��� xx��͝6[Ǉ�3r1�Cb����Ō�+��OA�s�a�>�� txKM�g4��Wd��a��/9��{�������p����]<���s��d	x��65A C��x�C��-�P�d6�o$@!#3�o&]�y3ܬ����W�o3������U�#�*�)���)��%�J�c�Y�b��	 *��($X�@�B��1��9��[%g�����.��-�
�l��@����`\.��A]n'���}D���[����Y��	�q<C`��̸�]
��B��D;����� �&����ncL}�d{�"Wd)��HK.�}o��L��πX�@4tm�1e��,7;Ԥq��e�����	H���((�9��û�!
!���8�x5utJ<l�k����H��q5��1)�O\H������\I����Y1�g8�{�i�q��j>=]�q����N��\M���a��,��Ϝޤ���|�<F1��07K��:a�	u��s)-�{�5>����΃��j[��{קx�-�	=�j"�x�P0U+�ݹʨ����/'�/� 6�%߲a����0h�~S�@�6ܚ�h��69Ya�4�~�e�w9Y���^��=�Cn0�H��R�$K-/n� �����@��X�"XЁ1���S� j��bYT���$o��N��H�Bw�wЅXt�V,�{P�f""j0'P�^��:u4���'3��i�<��{�wa>�~��K��.���>�"v�*�LĘ�#�|��Y���q뗴�2�Hw6|,�'��=�M{�1U>VU=c�F<L����fܤ�]ԯ{���E�mƕ�OE�Ѿ�gj3�Ŀ��q�Pʈ�AL�+�r��9�@@\�"�PR@	��"�!D �40�5,@
O�#�K�j!U8�՗[޲�iYE��j������
m��6�+���፥����ڱ&v�@J<�M�[^3e-#��Se4Ŵ"-��l4\�شD��v���9�4b.Yqu�m�6�Ѕ`�5Knm��'��(�8l/`���]��X�-l5�%�t���6��(����:���M�3,I�@a)c�̘4@�,�f��jU��6S9&���R��^$���\�%�@�v�qo���@$	B@��Q4l%���"�����x�x�����n�����&�䜗�D*X���� b2	i��[�m�2������4*^��5b`�@ssm�J��x1�^q��Z�ʊe(��:xf����!�����=)L�>b�/0�U�t���0��w;�K^�g���A�O�Kik�/�r4w�b��-´�2�w�)d���4�[v��t��Ȅ���l�>��O�Xh�5��2�����q���awC��nc'L1���n'��oG�1��'�<qh7.�u�� �u����(����&
�q8zJj:Dc$�^��8 ��,t��P��d�y�}dF
=��|�- �o3��S�q��c��翳�~r���#-�&��%� $�Ԗ���r�oL[�q�LtV��-�Ly��a���S��k�<���lDύ	~�b���z�W^��a�Z��\DHG�����±UUBxwr]�9u%	@���m,���<ό@��� 'qA QF4�[�Ζ|�l[�	�}m�4�4ů4od<���a���] ���w�.��}ޞ]߼�����>����]�)�����b�f��*�;dJ��[��.�v$��"�bp9�ie���kI��ߋ!��1�f<�y�`�����ږC�n��Y{�0W[��yL�	v[$���y�������jߪXt*:[�M��Z�#����SF33"A�� �"�Yd�������>w�|��'�0�/�����W��DX��P��t_�L<��[��g�ƃKw���ϲ�{�OW�\��r7/r�fi"`�"�����`��[���7%�F�*�j�R��x4��a8�c�;f�'�m�;Kd*���z���['ܳ����pZ�XPLBLb!�_ ��q0W[����N��&�8�����v;Ѱݗ��*��]O�����1�O9,:�}����/[nxFI۽��i�fk�-A>��}�ځ�މ}laMl�A�� KE0�����m�������-�S�Rvs�c��bD�DI���o�fo;�Ez�e��/�*�g%�舆 ��x��*����wt�q�2P]E9H,˳���鱍t��JIKV�E!��U�:ݛ�Mu6�l���[��DY�NI�w=����1�WT^��6@bCH�UץX���i<m��XE��8��u_>�5m�f�������s��pF%mÑܡ\6+���������^w=�����1>��dW��s���o>8�a�HN��<�8���W ��ZD��S%ӉxN���I�b	 yD�����	�[O.����� 0Z;�bؑC�5��R%���fz�g����A#hR�~�����i���O�ފ7e]*h|V-Z�g���C,�G�su{�ڈ�7���&Ǟi�"�>���)��'���5oM���5�(E������p�r���	19j+)�<�+�{���J>QUk�yUG�"�_f��Tn��Uh�T�T�ɧJrI;�B�&X�I�z�"��B@���B�3�LR#�*q�N*f!Ēd4��a""i(�"�)&�&&bI&� �`��%�&��`��d �Y$�X��Y&d��I$���p��,K2LC!�&	"d����"e�b
c\L��N1�Z(�&(&B��Y���b��Ѽ��_(��So�����ys��~>��6S3l�,�C3+s�~�_k�w*}��j�{ ����s�E�[y�[-bz��5F���]:�'K��e�rsbQ����]&�=н��(7ޯ�#$�eC�\\5�
3n`I<��>rOp��Ky���M�!s��`�ෞ�SI�~�ahoc�,xaO���٪�  ����͛�̙�߼�嗢}���߾^�ܷ|�]��a�ȌV)r�ZVԘ �6�%B�3�d\M��v� �2;@�! ��6ܯ9*�]�7M�1*1)Qȉ��Yyr7Ͼ���� 1$�[�,5�����j�:����Q=����9�<���_O�3~�}o�s�w�r�\5�Y�ܷe�k`O�OV<�`�s�Iy'"�jñ:�Uy���VJ�dxL�� ��Yd k �`{��,X��~}qzq�|��<�;��'˗%fo9�y�٥�I�"��&���G�����Jm ix�W���	(�A~�ּ��]�q��fE{��ʯ���,<[f��`n��s�y��ﭞ��������i��#QQN��0�����sXC*���v�f�6����� �6�P$w^.3���8��u�DT��4�rG����L�(�	È��.n�V�J�]�9�}{�ߝ�u�Yu#��]A����<*`��p��4��yܓ���|�:�B]a��LK"�A`�D���s&J�3�ʻ/%���|��HQ) &���+0j�(��J�k�R:԰��2�G��f6�*,r�nX�#�c���y>�w��\`��+-{�[oN�w��������S϶���v@� B���vëB�_= >�8aL�����m��-�Tp�`���s�Fh1ʍ�Z\��~{�w�!oC��`N�)�*�S��I���8}R�ٰ�@|���{h�۞�kG66�oO��>��� 
���J��l#t�;�#���V�B�]a�z�6��1�:xH�sr�n�.�Yν��^�g��M�������*�_=������a�d�(@wwn5J�nL�_��{�=n�>����/Z��i<i��ʃz�n����ܱA�W:`9�b$W�k���f���U7�r-���i��n:���A�t]˼Au���)(����awC��a�z]���=�ޱj#w��0�ViF|rۖ������G���=C�����Z4���\5���
�����O�2`  C"L��
 ���ܜ��R8Ls2��'�M:6��<�94���A���,�'�}ɯva����Ѧ���\�m��0�1�*����Q�xG8Q��0��	H��q�A0ȡ�K�� ��L 2t瀸`p�$P����:Ȇf(�I @�#�D3���*`�(�\ a�q��&v�"�.	E�"`���B )�*��VZ�U�`A�X�-�P��E�,*� !�� g �r��"e &R"i� #�"$"�@P�H�Fq(
@EBCY��; LY�Ñ���d��%�"i���~�˟nH{@P�"y� �1	��IP4�&�Y�Uat���APf���E)T(R�TR�`*hB�W��0ёʳ��d߀���Yq��7ۣ��<����`������	�h��q��NG��J��#S,��F��3'�w23/d0���.I�3s,'-A��5r��p��9�D�g� �z9!��'�&rp���}KE_8)��ߟo����ә�L���~�&�	�w��|׊�g7����@Gǳ���vS��E�������L��Sܠ �#�P�$�E?A�D$�4	�L�=���ߣ�;W�v��3^'��� �vƠ=xy�@TP����� � � =G-Dx?�x��2��t(Ni��I���z��6��AԠ��E@Fn�[�ʪ����x��N������3$P}��4x�Sg�֟%�}�����y�h�v?��VR�1�9��L�+�$���=�`���NI�:����#��3 �߇<�S��c��L+�=rp�����>����k�c�3l������L���{/��������:��N��Rh3��{�C83 ޾9�I�E$� �C�`��!
��6Vr��@bV D�caA
��*
�T1	@ЍHP�I�� C�	�%�	eA
 �Aa� e!�)B�ZV��(A�T�@D�TA�@BYQ�` V	XahbX�a���fI8)��)0�ұ P!0�@4��"��V
A1 bE�h6���iM��@�<�3�c��b Òl��u�O�sC�z��=>��6F��z��MO����u8�#� �	�r@�<�����!�uu���<�����0=���N+�˰����"R�g��.]'q߫Ф'���f���N~�����\��>����9	%��z=~�A���>��/W�G7�>!�G��%���=�?����}f.���m�{�0%p�$�h�����������(���������������������)�����������������������X
�������J��a�(JI)(���a��Xh
JJ))(i(bJJJJR�����������)ihfJJJJJ ��������i)&)) �����@����J!��i
JJH��H���������JYe������I(����(JI��d�(��bH�������JJ��i(i)&))(i(bJ�$��I
H��d�������ZJJZ���JZJZJJJZ)
JJJZJJ
B������������������b������)(i)(����ib�����JH������i)h��"F�!�JJ��b"d�(i(i(hi"J(d��������J���������������������"$����) ��hh�)(i)i(ihhh�JJZJJ�JJZ������JH��!��))(bJ�������$��(������d�(i(i(ii"J))&JZJJH�������e�(bJJ"JJ���!��(h��(bJJJJJ
JH��!������a�)`$�(�����I���!��b���JZJJ$�f(&JJH�!������������	i(h��"��������������hh
JH�JJJJZ))(i"ZJJZH��ZH������a��$���ibJJ��"!��i(i)"J))(hhbZJ���)(��!�����(�����i(ii(h��hi)ii(bJH�H���!��(i)(���i(i)(i"Z)"JH�������H������!��(���bH���!����� (hbR�����Y����a���"��!�������))(hi(h	��������$�)"�"i� �������"
b���&���&�
H�����


���
ZJH	�`<��� ��NXu� �
h���x���w�	�|���A�;SFq4~������>�?�����Ò�<���d^��Ӱ��ϬQ���z2^�y,/|N����6��;�|W�#�G�6���D���K�Oj���24L�x+�Ð��ǵx~�x����� ��t��Me<	� %@�BzT��}j}'Y��f�I���j�)��aǍ�G4��C��=X`z{_��C�'z�v�Y�������0����k쁰��FB��a���=0�@ѡ֘G�c��@���?t��]�>�;L( #��!����t}v	$ ��&��C�5ZZY0f'��?T�]�0
�,��'c�Lyq�F�����l�~��l>>>�6E6�[u(���ds!����-H���$�	d'��p�	���u78�� 7Sq��}�$d�G�>�>|�x(C���8M���o���� 1� ff;� s*�ta&0	��*�	2�c
��#���q�Á���Alt	� � ��T��@� >�A�H�ק��>IQ��͙�mS�!���Lg���K����x'g�m��̛�����h�'�'� O:}����{͗ ˯�#������=��%������L�U|C0��6��h?��~)��D�6�N��
�3<�{���Pw 9�ı y�#����|����T��㢦��rnn����O���:����#���j�#��$6���G
�0>`8��PuV �H �#9��?��<}�_�<^8�&�Ze�8!�6(�/Bv)����I�pOp��!���v��y���z��	0���qjp �댃�8n<������i����`��jfh;�_����U v��~=�Fx35�<�>p�As�N`��[����r}���`e<w2��8�C@ɧ\�L��HM����7�>����#�М�`2^J�_@Jt������1�������M�	�M������ ����"y<�:�������B�/��������U�UA�1�` �J�)����0}!�"�	�L��:x.�s4=G���@ G����N�z�"j'a�<pǎg�}k��\�����^c�m��=ɦ�����. w��v|�VA�xiNx<���l�v|ۺ	}5I���}�R��_���"�(H}M�W 