BZh91AY&SY��\a߀ryg����������`�^ /�  �  �  �<        `  c}�(RR��Bp�GhH�b5B��B�S���EV�QAչr�4�h���E:�\P������eƍ
:&u�QG7N�=��|�.�(���:6tQ��CF�9�qE�M=o,Q@>�@}o�PѢ�[�(P�p�*fӔ(��[�(�(��� ��t�t��qES�9*��v^(Ѡ9�qJ(�7[� ��O��(�Ү� S易   ���              i�)R�D0�F�b`F hi���R#*�M6���&���0�`�M4�eI)T= �  4 4   Jz"�����  hL!�aD��h��hM2'�a��DzF�2m1������Q���L�FF!�C �#& ѐdn#ˬy�=����w3x� �H�Ј�!�O�V�R袢�%��?���~��`�I�y?��-������o���ƭ����kU�s�?��f�q�mKp	�r�uM�}4�\M��e�K �$�z� a�K6]���2	�y$�x�D��I�oÏm���̠g�a֗.�����USb2I�U>��c��������	÷i$`:$ޑAUP~��Ar:P������ߛ�J������FI�'R_I�K����=</l�Xg��H���و�� ���$����Th�����}��ux�r��>�\�E{<QF�,Q]�k�r��+Ɗ4RW5�+Ǌ(�W5���wy\�+���ww��ww}]�k���W4Q^�]�w��r�������;���Qd��﫚(���h��S������i��s\�Q�W+�=�������Q�QF�+�(�E�N�����\�PQF�,W+�(�+����4����s\�W�W5�4W�5��x����k����}��k��
(�ww���ݮQ\�+���t�k�(�E�Q��<�\�\�\��r�k��s\�W9������W5��s\�W��r�]����}��s\������r�^9]�{\�+��r��Ww{\wwur��W5��r��E{���ww}�Q��+��u����x�\�h�h��k�����+ۼ�ww}��5��h+��r��W)�R�5�4QF�]�z�w����]ww}�k��r�N���+��ת(�+�)+��;����k��r�4R�����8 �s��9u.����9u�r�N�y�����+���_�s]w����]5���u�(�J�r�W5���\�y\�/��r�^���s]5�5��r�\�����w��5��^<Ww���N��+�����}�|���_+��r��W]�s׍�r���\��r�]��(�F�J��5�(�r��W,Q\�+�z�r�z�]w����us\�PW(�)5��򹢹�w{]����\�+�(�\�S�����Mr�e_;�+�����]5����ww}�Ww�滼�W���\�J�򹢹N������r�Wr��(����\�k�뼮h�k�+��}+��s\Ӽ��+�(�k���+����;��ez�Z��\߲�~<߸���`��=x�x��!��y�9\�k��\�WMr�\]�r�r��Ww��%r�W+���\�\���r����\�+��;��p�W5ҹ���s\�k�=W���sF��W+��W
�\�w��r�wy�RW��h�\�w��sEr�r�W5��W+��r�wy^�5��\�k��^9\�k�s\��W5��G+��r���ҹ�����|�
�~?�}�k����s\��r�K��J滻�ﺹ\�]�Q���}�Ww��\�i+��\�k����|�]�k��\�\�}���^w���u�k�k�����~W(�Fżk�ܷ,X���yr]�|�  �S
L ^P^~�\;+7/���s�8M&g\.F���~'gnZg�u��ÙL-w�F�����U>M�~�Qn��Kkd������`8��
$0L:a�^�^�3�O�0jqU�⊵�N\�I���5sYn�Z0�jbn��c��i�����T�}8}1E�ba���1��r.�عQS�!�q�L≇{�9�ڹ3�� ���aU���"rnM�\ٵ8���ǒ�]\ø�xy�/":!��#(U<����䩘�2f���B<�|J����#%�M���*���zx�-�����F���(�te�X���a%B�oo9~��-�ʞ=
R��U	��FH��W	<�]R�pB��
uue���Ӫ4TK��r�b�fJǥ*�c�
��rD�I�w ����엷k���6^�*Uw�*I���IG��jjfh���pe�S��9T\��o)ŧ�%�C��Ȍ��CYq���E�eU�n`X0.��'���Q4LF;���F	12Ü�s!L�̛��z3A;P�{�&����R��>`p��rIw����w(�� ������N"��*���DKڸ&���zLZ�Q�SX�ӺɌ�R��9���a<�͕v�\�ȜxOt�K @�73�R����r`�ˢ�pP��7YU��1YH>Z� ݜ�����UQ���J|�i��E���WrZ�(���!��Ѓ1oF%��m,�n�= p�*�3���Ũ1c �sp^.�T!oT��\�C(�"�s�3+*.���n�*.q�Q�p_$Sٌ9�o.H)3 D=�"���Ww"�%EDX�ɷ��r��]NNFX�
�E��j���_��h˓�՘��)8�.D���f$0`��t	��T	W�F!0*X�9PC�P�����aYy�Q�Sg(��|��jH �e���4��[��Me#Lb�j�Zʘ����
����j��4�-c<�m�ҥ/���̇����*p�.Ӿc��^���&-H��^!��B��]Ne��p����*�m9�c2�(E(y�B�Y(	�l��*�"1��%�(ò�9�yo5p��2�
*r	��3v��h�9*��TF@���U��I��#)eG�[�1��SU3����`:�r�d]�@����S>�ARp��1�҅�Q�ʛʸ��q�U�U�[��u��/*�E\�%�V�V���r"�]ز�Y���/��s"�&���R��w�'�O�!��.���/tU
��Ur�	��Y8��"k�Te�s�dR�G*d���9T�L�˸��0�8�=b��x���J!.$�K��⻷s9P��6m�/1os)�Q91��T�&��oy3youu&.�؁Ss!*�P�A<:�9��=�9{*NT�x('��
VLTc���a8�[�<�S~�SF�j�ֲ�]�9�1��E�Sj	���^T��dM�F,Շ�r1�T��
��|2�J��i�b'"	UFU�3Yr��R\<�e��NfD�y�YQ0&aD�����yn�`QyT�\���rdU���j�J����o%�$)�BB*rr��$*�B�Ș�5�]�^�6����]`F�|ˢ�!�n�)�)��9��m�.���v�ə��6 �$1ޭ���:x�PAX*��!Mc"�U�
x�X�X&�L)s5������f�20�yv�%T��=ϡ�`�����?�?c��㒧w*m�7*Z�*�0�J�  �`� S.�6e��&J	v��  �+u� V��	rX �HU܀
�7@�` �X*  �%�J�@eeLA��
�.�p))  $D���b�Xبa�D�ܕ6�PKD7wkD$Z`K�Y4@� "�]���
I X�Ar�������
a[��	���� � ������(,���H6f�!7wK�A{���2�!��*@�AHU�@��W.��+r�kwA��}�<�g�
���%�Χ������ki�����a�,HS�7i�>�M�u��<G��������И0ΦS��p����ۅ`�'
!��������<�2|�2r�bx�����bO����4>�cRkh��es.R�7E�dh�q#.�R����]hf���0�*��݀6�i�[�mhT����a!Cl�p2c-Pm�v*50a.u����H���KQ�Yԩ%�����������&өf���6�����څ������8R�":�M����f���f��v�)
ؖWM0� .�+.��7���]�LU!�m�
7��
��T��L��35L$ԍ�6��Df�Tݪ&z;CK�:ʳ��v.�vu�4�9��Kʹumq6V�(�p؛Z�6�Y��6p!73�lʪ:ݥ����5e��v9b�ΉXl5�iRl]��X!d`[�
�k4#��պ]�h��iB�h�GCBꄢr���F�jS[�]��D"ͬR�5
�.İPa��;-d�Қc^���lZ��)ͬ�?���{*�e�ڒ���M̐�[z]b4+�8�if��*0�uz�I�˭K`9�Ìۥ�6�]LRځ��Q f�I�9BP�ʱZͮ�[��eu+1c�3�;����V�(bd�wа��#
��%R�&�h�͎��JD�����f�5b7#�t�
�Y���L;Z��ղY2����8���a!+)V.溛�Gjl^!.��׼��b3.nVBkq��H�.CI4s� �P�-�gM�*Κ�6[�m�[��!��ek�3�&�a�]	"˱����2ш���/]N�f�����9lL^mbE�֔GYk�N��D��g���3u`����D�m4����ٱh�s��Xg(�.ͭd��di��ԕLd �����r��:JJ���PКX"b)�^G�RR&P K)�ֹ��R�����,1]��b�I:R�A�.�K�0òvhv�kt�q�	CXa5in��6q!�qf��b*)��M#u�`��7�v��b��1��X �mtr�L4n�qs���ZS\V���J8�+�GZ����h�Vm���A���D�G2i�!ZՆ\�l�CdB��a�S��J�����Fպ\�15��掠�\3Z�h	v�6t�+,js�W��;J6�մM�R:�]2��n��R�����I���Ml�S��`_������&0x��4VY��L��~#����[L������,8��P�����w�]]u*��������=&��^с��(;�n��ky��n��vIGuR��=pe�m����I8P�����;=_>N�=k�K���<gy'(�Ĭ�L��|���i�T��<�+��'��<ӗ<���P��S2>��d��B)$���GԜ!8�V��G�~<E�׉�>C�m+��VF���I"�$� ����<�N=�o��}�Wԏr+=!	'���K{凄<�#�N^ӏi԰�E9��Y�l�o<�p�4�Y��/#�B�y��������W<|H ��OeoK�D+t�������ޢya:N��)���Zo'��!e��k�C��u���aǎG�Hb&V��AT����-��z��	���R�N��[���Fac�7�r|g���ޕ�'�@���JL�e�*x3F��ye�G�ӷΕ�:�+e7��|����)� �sM(��9�Ng� yq�.�$[��c�䇺�+DŠ�L���'��q"�fQzx�,P�P�i�J@˻��R�����d(���D�U'0��W�f�����R��{�w��2��GΟ��N�_9ٞ�ʯ��4�1���IeC�`�LPyF]8�n����!�6F>D��AD8<XUH�y�p����ʂbN:����wLf>fL�N�Y��޾=���
ǼMOn{wߔ;���d>=͜y���O;�'T>���o����/"�S^#$A	1x�E��渶��cW�Н����_�;�{��}�zf�-�ڗN�r�2��9��#
IWI��1[���?��@#�A�mx���wbM�(� �*D˔�9�aDť$=�h�]���f�:�wu�wZy��6Ի�{�᧿ae�k-��OwZ�_����N�k��<Aq/�E���;}��r��DR:ޛ$���G��|���/��g�cُ.��oBWNՠ{w�*Ϫ����=r#¶w���~�I�%н�N�K�C����T��a=]:���2|�Wϯ)�=�R����)*ac
�o�&�qҭ �ʆD�c@2�U���1oՅ��0�����h�B�A"Vt ���Ǔ� |���%�y ^���i���N��{�ϓ�u�x�{@��ӹ@��x�}=�n�2OCN�g����t��^�x�U�ԲC
E�cGLi//�*g ����<B|'
=�C<W�3B�M;�C8���c���y�>;��U@�@b�I$���-�YS���gR��$�׾䟙�7��EA�l��&� VH���K�V��HD�
B7f�)D V��@E��eF��~����-��~J�����i���ɲ�� )B�5e@X� �K�&�P#$�����MUZ ٳe�@]���(`1��v��I�<yg����Ä>�d�}=��v�ٵH�Q��\h�gkF��PF�a)������V��sX�&�-̔�K,��W���i�eI�m
�f斚���K�9pZ������sikX0���m��Y�9�2Ie��WĎ�����,��ծ�[Yf��7%�86�4�e@��G� l<fɛk�h�(WH]��FSF�Yն��5$��ڥ(�ۉ�b��6�]�]��&j�lu5؎1(̻����; ]M �Q`� ��+"����$�UJ�I�q���Y+�t	����H_�Q{6N~o�NR���{~U`�P�x���fCK�iN�\��x��� �6'!�{N�:�lp�ܶ��h4����2C6�	�E�"���Mm����Cj��{�YIJ���	������m,7���q�����v�ث3�擌I�i�oW�65�����8--�ٷ�b�2�*I'��a��0� 3:O��ty��Ś9=F�\A�L'>*=K����I1z��z�n�ê���ڙ���Ӷ["}~�=F��7{;�ܙGar�SY�̛�������00���@���6���׻7|)z�Y�	qq�t���vx	����x�`��l�v|ޡ�A@n\s�cU�:��Q�p������=Kim�z݀M��^hj�X�>U�A�׶(�B��r#<�e�7��ס��-�u���@�60u0&���ID�@w��<;�����\c�v��,)��(u�#�Lެ;s���OU�I�}y��]�߽|Ͻo� H(h���J=�u�18����B�^�'}y^NPH�@Xٹ����6Ź\Q�Ќ�c9-4���uY�QJ�)����Qz[�X9ۋN�.67m�:��N��B(������A��۸V��}���M�b���f��٧t�m�� T��<�p���@1*"!@w��Z��]���T��#��Rv���>z���t��O��H9�.˾�6f��nߜ��yO@my�L�څ�n���ߟ'k�KӲvgi�r�.v/�"���00�څ�ja�v+���:�%>_#�c/�K��,��1����7���(��^��Ѱm������ۑ�fDpY��6���I�7�5���a�l�}=3z���u���<�B��lC���Z�c&axd�!⦜n�3F��@[��*Awx0���� :!�J"h�XjѺ���m8	�����k *���yT�k��>y�>��NW�:����Y���a�" D%��\I.H'b�$٩�]Pp�$�3�^@�HԒ�B"e�í�SFʍ��E���]|�S�㊵H�f-	M�2���M�[��ɻLh͘MH��
ő�X|��|o<��L�A���l�&�P�C����f��kʦ����[y�z����y/�E�R'���*��������z���?��]�zG��>.b��2��U��W/����o���oT1��D$ a)a�UoO�L6�����@n���0��� O��
�-��
fy�P�;�k��$�-2$�7������z���2o{m�ր3�!��X`''��l��t�R΍g�S��v�ǚ9��2�RIc�Qq�`T��J�ȩJ�rEc��|DǞq����^E�xǧ�.��|�����jh���X^��|����#�q��)\�]�W�����f
��� �r��=��D�P�km������M��Q�C&&=P�|&2���73J�p��W�N�2 � H����"3};�ЁD��Zb���A$YHHV��c��ݏF b`�x�!����G���a�psro�@�3/-!AI(1a;�xr��3BO
����-�{.y���!��_	@���nm1�fً ���l[X�@!%^	�W��ǡ��9��&���"���7|϶rO��������7{;�
��a�U����	�q�0Xҡ�'�S
%��*Ζ�>n�\T$8�َ�1� pn��a6�#H�:Y�k�����Zm�{�~oV����d�e��F�]��uU"�s}�Ȁ"!�DC�`֯�:2�vK�8�&�r:�HJ�V�ɺ�*B�dW�RK4X2=Q��L�����-��l�ܺ �]�`��+��xxv� � �h
���rA��E��v��8���ڰ���=�f[ �,�-Z�l���N1-��>j��{���s�kDȤ�	���i��v!��<܁�!2��!J�z�@��ɺ	�B�2m�l��k�@�C�i�[k��Gb�g>���=?~��M����qPZ:�G�%<*oc�p�1~f�""t�cd9�4�\HE:|H��[_e��||{��[Vũ�3��i' <Z��#�%<��D4�lu����$�;��a�H˵�Ӄ����'��ǟ|���Yanh��GHm�m������n�`��m�HZ�5(;8�FD���5�N� ��,�v�D4� q�"F�k>BxsE�^e)!��f.L��/�^y~�Not�����,�o�+c���,�&Wd)��l�Y#���2��5��Ѳ����$�=�]s��[P5s�D�"D@J�K�<»�2�(���`�wq��1�����7SY����qp�ɲ0E�n6`nY�t�I$��O#ȼ���a��j����cZc\j��E�!��
b���΄$@p�i}�)n�
��2�7��KYo�q���Q�z��-�t�U�ql��!��v}>�ܻ�{\l����<$�]�ڴ�@�l�����q�<@�G=nr���ya�X�0��3�n�<	"-���q0U�q��j,6�]��O1ʧH���#���L%�G��W$0$�흳�i'�����y� Z�8c�H�w��Y��=D��r�.Ӱ�)8^sݓ�5J^�����l"?sҟd����l��7\���4ណ�84���xP�ç��J!� AcP@ye�`X%4x{�dw�+-�Q��Z��ԷlX���Z�n&�,4��f�^�͓F�2��N�{�e=D��-k�;Q��q�SD;��V4D��%�p�,�ϗ�����G�{!�����l'��p'�5��0�c̀x�,4�[-�D�v�$��|�y�'w"W�:��*bS�0�,V�",hj�� �(�""�I�Y��H���P
 j�%���c߳���a.�.����̜���Nyȫ�4aux��˼y�q��<A�X�G��SQ �G�&_�DE;x���������D�eR����3ըY�������V�=l�獩��1�{'k30`^#�3>|��>�G��zjd)����<�zC�xI���/q�r#U�ٿ>���x��� B@�E颀�Q) ��D(DL2��،7X�X��[�4���b�ˇU��`T.xMn���Z�U��3s��d����-M�b�-�0(�s�7{�J..�K7����R�#�mV�m�d��\镶�%)c�SX�f9RR�s�
JbQ5-0͘���M�h�at�Y��K��1�YA�q]fk R��L�VjԤ�&(9�k3M5�Wl�ji��ݳdv�ڐ��\SB�n�e]��6��!����]��5�7e�:Ϝp?G���c��
�~�}y���Ơ��FŢ//�fڸ�@B��y{��pҁ�H�b4KkCCV��2!y�G�6�E	5�@�o�ᣇ��nބ���1��îK�f($����ws�O��K����&���1�XD��\2�Ø�+�'Ha��-$^�� �ǘ�ܘH�8q˷�-���'��� @�v�Aӹ1s$�����i��;�>��}��%����}�X?�D"9em�/:��}ju&Kh�����e�-l���4m�і�Vt���k��<��Z�6��=L#����+�A�T�u��64�E���_\K��ɠ�c[�����
\%X�����ȄnV���c@��7J,�GЃw2���OH�N�p��h��@�Ia'���.h�$0��O�_�s�Mϝ��N� ��i+�L��q!��6ǋQ֢���s )����Η��gh;�я �2�}�NYqr�v֖�'|����y�qn����m��a�xŘ	 �E�v��t��Ӑ�[����	a`-c��k^�@��8��%�I�-��k�ǅ3wT�� @���!8�S��r��g|�>�3���9�߷�$�5V� J�OIv!?Se�,�Z4]�WMl	�X�\��jBb�yt|�
�G͋:����ٕX�ۢ�\$��i� W�Vx@�������q��b�ǚ�y$�,������O%<�`j��H�x�W��<9 ޤ8�j;�"fe����8ˆP(��<�l���{�)ϟ}}$�8)�%����Ԋ̙(�-,s���O��'�#�D�އZ��T	#K@���=��4D?v��d��S�8�un��)gW�yl�9{��}�vF�$�=��YF@	�v�ڝc,zH��̫�x���b��3X4b�S�Hx�h�1�F�[&�4	#����U�6.Wb�3`ɵ�]�in4t�l>o�'���ƀ����Kil���<T���x���{�Yv�F>�b��И�4i��t�B��OW�_�m}�����m����ZXAh1d�v��tD�4wA0Uk�a��j��A���O fS>���,8�#�Y�m�qh���� PL���$��nu�v]�_�o���;�>��~y}
�VH�>�<�]�7��5n+�L�Q�d)����Z~���/��FL٤���[.¤�h�V��x�;l4bb1�;F��y���$ܨ����Q�Y��`��.�:Ũl5�"�h�YJm�QM��OM��@��Zƅ��l��<�L����F (p��P�8.��-��4V���$��eW�zz+�>�â��:�M�����Z��gc��k�rz�k�,���'�@�o�$���B�d	q��=�����[,�(gTeSϔ4m-�ػm�;Oro
CN@M<�|yD��,���Ժ��N���'\By��_޻u�yp�XQW�;�y���>����>{uj�L\��7;V�M<�_��{�/�(�v����ө]��M�M�w��Z�\Pכ:�>�F<n=����5�,|�.0��k�T��fG���MZ0�O����Y�?�h-To2p(�P���{�s
�^PWot��Z��OK�� I8�X�����$$�BBE�PX�j)#RX���V�	%5cTkb��dD� AKDqd�%���������0�U�i���'Jm"����9w{ص�V�qv��A$�O�2đ��
#�H=�fx�,�}��,�Ƙ�v`0�Ӑ&���F�����Af�/v���04���6�)����}^��߂��I��72��p!�"
QC�
:l�᰺̍��m �$�ѷ�[����$���AXņO��,��FZX6��e��@Hb2�XQ����R�.|����׽ɱ�\㯻�O�h� �b�]v35�%V�L$GR˥���Ԑt�'Vj�$�h"�c��:"M]q�l8�1�ݤ�r��+PvVG���x_�|�[<�u�Ӹ���)�)o<�aΛf ��$B�i��E�ů4od8��	ZY���w��0�f�]$�

N`8$��!��1�	����IWyķ��OA�`��ଧ��D8M)�=x�w%�ǌ���0Kw!GK= �{���1l�Z	"�O�y������ĊD0Q+��9]���9��ެ����4�a�:�����h��a	�$ĬNoUM �����1~�5L���}U�	��7
a�x�{���˶����l�5U�,��-��'��H�2h:l�i��W<�sr�if�;��]�v�n󁘇��0�s"�WWQ�oI��.�^G������[+8�J�R��mɗ�������B��d����!�S��K\�Z[����g��=����� ��wd�9��ÓY�~1" �Y�Ebo��FJ�ˬ��]�z�'/��ߝ��u�Pb��,":����-]Q�vu�Q�l��gK��0�	d�Yl���m��塥d�x;�@��H�qh�[˶���l��o���w���aL���Ѧo�F�*֛ O�1�f�4����xK�Kq��U>}����g{tQ�E�mќq�����B�:��i�Kip=۪ h���y�ɧ��8[�n�[NF�sc�[����a64�#H�����t�PS��K�w�g��K23q�6۶;�w�i�$�-���q2Q�R`Pt�E��es�'���]����Ø/��<�c8Ip��N%�rG�Y޷���@�M��7s�$��@wpDJM��wKd��o�h��/���@�I����&ߙCS�0h�u�<h�m8{H=���%��{�X{�?n�Ȭȷ���h �3n���R8�6CiY��ϱ�{��;m��̧��z�%��X����cþ�@��y@�p�~?s�Ķ�GX)��[�?!$��-'L�!�;���t�T�4���46>���3TZၫ�%F�@%R���9���֌��y�s��C����2"�\( �m��9��qDA Z� j��9�@OfT�ɓ�f|��_�������Uqރ���(�E��".��O�Bj]H� �&0��b�=g�x��} ������15�h�ߜ�]�e)�p���0�C=qV�U�b���V��kB�H<F{�p�t�ˇ9��=��Q7q�=<>E�DdA�OT}H�0�TT�:�B�<�?/�K�˺;�[�w�ڪŌ�#)IB�Ich�-�0�5h!T"���@ ���\��V��V#( 5hB" �#!ifD�g�vV�qԊEl�<�[�-M[JGA���RPvn�7G7
E����-3����7$E�	VV\�.ɳZ�Ij�n7k�[��됆���a,�v�)(3]����V�ͬ�e��� �l��I�h3XZgZm�c+*kF�^h��i�v�u��tԶR��B�eV��uVQX�4-�(ݷ*�.����v��t��m76��V;��d�B�u�9ҩS)FX��Rc̣X!�RB@$�FBTQ��X��%o˕x�D`��-��Z�Ajq�B�9 I	"B����뼿$jA�%�%���/t�E��dfڬ�8����e�ֈ�)�3V�e����(Z�Yc;e�#4)ayd�%ƚmj��M�l�l�x85I��?���ӟ}^$i��?6x�_����M1��b�ǡL9��o��q7�i�Z����x,���pX$�-f}9�Fw�b�a���eQ[䜒]e���'Ht��|h��ao�L �nn�x�Cg�E<��¡]�a� 9�E6f���j#��mu� ��<`�_���~yY�0�� C�D3���C�v$�L��N���sߎ>��*~��@��egK�<t��<@�SPP.%C��[Y����`  �/DK0��Y��ּ ��r4�0��l��*9��F�ܨ����)g�ϖ�锷�t�Jm�/�w��ϡ����#�·��!����Hܗ��gh��.���������{v�|!0�g���]�U���a�j�v���	n"H�	��Ʌ�u���O�-�˗,8Ѱ��{������)�b��Kx���@5�4�.���� ��.�ے{�����>|���<�>�7�>$$���E�(���Z5c��v5\�4)�sWg\�l�%�k
r�0��踃cjk��	�w�w�c�K�z��y��K�c���AH�� �yR�K	c��3Y}=���F"[���e��Ϝ1�v/�_�Q �6pq�.%�#-k�)�������&Q�a�ir�pç�ϗ�;�Yt�U�;���vh�Z�}b*qXh��O�	�j�g�<�?<ߓIm0�p7�ai�iZh���à�rkɔp�����on��Q.'���u��D����[�����k�8w,{3�
�� ��=�X#��D�}Ɗ`wv��1�;�i��eˌI���6��T�1ݶ۳r^���.�7"��_9$��&�<���a�� �j:r�R���0a4���TuГ\w^��A�Lua�e�i.�-`�������_�MJkǎ��Xʡ>,�kb��B1G(�������<{��<���n3�?_Ki���>,� ��ߝ����0n��:Z��E�Y�ky٧�`-7^_w��ߵ$I @+vlы@�����*��L��d�n"���X�-�@�%rb]������+����g(���vG����gĕ̈��ej�[ը`\�y�S/!� q���6H,a{�٧@ Ao<�{�y�Kqkia%6�[�M�0@Px�G�@)vE�7������1��$�{vۀ��ܪ��c׭��/: <�a��v\	�@#w��eu��"��@Ò���\<�$
\���
l�Ƌi�F���D��t�1���Ⱦ份ꣅA��b8Y��9�K�=��a�l��[~ �������Чk�j�x�U
�9YV���WD��1U/���V�UO��5sc���:4|�+�x�r&�;�e@1RiNg�ڢ\�b�;>�{ٵ��j-ըyQ@�����<���mX7:��-e���E�7Y<��Q�fnc <��yx��%����F/��IP��JQ�(Ǻ��]������@؃P`��XذQIF4$d4��-%�F�Q��a2j�h��
66d���jDQBȩh*�� TBF̐,z���� Hc�z}���4��������	ގ\���b����y@x�&t;	۔�!��}��X�P��Z�E��?	���@�:�u^� �:�3����XV����T�A��" %��	ʈ� ^fY���;�#Dod	�`v�; 5�}�g�i���h
�<�!N�|]�6���yi�k,�4�@�$��$�3�ws�hP�x���.�.��O��(�� @�*��-T�s4����.z�ᅸ��ZI���2:�+,�J�0�	b�ɌYM�*����mu"˩w6V|�����yS<UȞ8��c`;'�{�"$V�Ű�oeD�KAv4�zy>��������˳Ȍ�f�̗��wN]�!�O�G���x�W��O�\o���(�R�4FLW*����'��`�������2��0h�%_8�p��V�h�33"
F�;õ��$j���<������������Q��a�q<ũ��pR
��>版��S��8��wͅ��<��mTCq�R=ʾy`.��VY{���ș����̴S�/����4�<A��-֨>`@Ƅ��w�<X ���]Q G�ZŎ���Y��
b&A�i+lv��<�j���x` �N!��$A�ye�ϗ�$��>�p'KaF�ЛDZ�b �K<N�;Hmc'�=�L\�}��>��W��{���a��1��5�f:t��"�ܥ�����4
� �U�/�m�L
&q�5YqAc��Sm���E�2iaH,E�TΗA�j��j�]�һ�0NJP��khH�z8��=�n&�"�V�t\/m���Lm�0\��2�a��j,�EQF����c�(2�|�����ʪ5n��7��a��4����Amr���QlI��'�@�3����.���$E/�I��V���k�\
��Tܘu�6�@��ka���A����$�ލ	���ecA��9�˹M�TŃ�=i�>��i �n���je*�o8�nP�ΘY��V�t�������v�a����1o�X�+�<�b��-	�n�j2�2 $R�J+���dr��j���y	��g>�~a��^vM�0�	э�x,*��"�l�x�+�L��L��T���"I1%��Yu�s�yqNF�<��<ɗ���-r�~��4
��xu����8x��P�f��a���  �-UŁ�>gTX>|��E��O	��2�9*e�.@��xoe�����hs��V�V�"�R�6��X֬f."-d5k"j�B#	��b\ơ��/�~sf|��^�6���G�:�1&���"�Ϫ��AVX��-b�żyzޝ�T�<P�u��`��"��!1�s�>�f�迯��ČY�>���������旧�["`��Suo"G�>'��&2�L\?��K�
���J��dF]<Ґ���ǅ*�<_��X���tiW��e�I�j�D�^w:�U�U��I�#6--k�@T�C@Z֫�4��&.�ы�"]�]XP�LX@L�"�����6s�7��
��!�[1C-�U�*����H�l��9�R:�b�#��ɰ<Ie�ٍ�]Q⁊�A�˴�n�v�R.6�E��2,.���I1L�ֶ�Ť�M��-6m$td&��iH��ck��a�3s�K�M���L������P͘�4͸��3��B�mca�њL����\�WQ���i�Ƽ����[�2kr�EJ&[�f3em��.q���h��{ߏ��bp ���;${��E�}�_���\�*ne��䶁�L B"H�&���DJf�%I���3L`�Vj8f�eJ�"��dsP�荹�4)OXzs�cw"c1���S]�-.�'�Z$�d��I���6��0���=}p�K�`@�\���i�ژI`Zi�+_�@�.�4�~~|��{�����`���S�O�*�c̤�o ��n'��$�F����2	S��������3�	n ���qϛX�+�ī�ՋL�@Q0�c��8)���9����3�TDC�+( �.˽}��������>M�c��v��'�M��i=��,3t�颪зp����3��O t��8h�S�[��- aL�\: �
"κ���m��3�o$������w\DKx�>-g�<�}qM�lel@�:睥_���,���f�$D�q�{�3 �6�VT��E�)"؆]��U�ˣ�[��le�ʜ��Z�τo><��e'K3� ��p'�,/�Q�&
�q X��4ۼ�+zN{WS�U�o��z�}�$�! ;�$!g���v�t�I�Ѣ}��!*��ZL�����-&�b���$4�M�9t#��e�i:N*1�g�䓓� ��ȫ�Gx	B/ ��(���a����ݶ��j`�dނ&���e�ّں�����xv��#N�ݜ�vw�;(Ъ����&��S�~_'/� K��^�:}�H�YծЫ�eה���0���d4q�\Kalf [f��R�t�0���J��K���_�?<����;�벉Y��6d�D;V��7������`��1�on��`�ga
8p��Um[�Bӻ ��Ir��O7.��"·3�n ǁM����B2&""
p��O�C�a%k�vYv>��f֖CKI�y]<�j<Ũ��t�5� Ck�O�a�hL�����*T�3��0~����|��|�ߟ>}�=� w�c\h�@�R�^"�� kB���ik��ǣ��0��gŀ>X�m먖:�(�a�����nm��`���]��"%�L��n^��%�>���7��u>w~w���B��҉n�V�ۘJp������.�-j�t�b�%qXR#��v�BA=�y�v6��n��b"ds���s��^OwÃ�_<���m3����h�N��0�cͱn2t� kI0����cbSx���~�����1�#��\QR��8-����Q�w��O1�#��s^Z�V�.Ү���>!�4h ���]{"�7��Ȗ���̋�g��
�����^t�t�+y�����q ���s��M�ݳ�q�?|_�~=����H�x=��v������X ͢J�WU>͓��+��FE�T�f� ��^xڨ"nǯ2L*w�5�j��uK��)��<Y˗�ɚ57o�
�����P⤡��]R�'(�^���Q��b�/R����[��O�U�UdЁ5�&=����ҵE����/)��ro�8ʒ�
c��y)��0/�4����jz����o�M���9S�{��CĀ�,� �y��0�y��y~�?#�6�lQŻ��Ki|�@�=�Њ�\��s�ۖ��e�c
�Zw�|�9�V@�u�o��-�����i#M�^~y�4&�@i�e���6���%p�f���A6��p��vR,{ELV1U�0�0J��.��[�tIM��p%���N�@���H7�Fx�GH� ��~��clt��CDj�S�䗒uu��מ��hB��f?s8$�>7�5�_]��8q""D@��UW-ƈ��ڜ�p��dm���λ�c�E0�m��Kn�m��e����e��ɜ&��@|���1�9Y}j��,<eә-�5O<�`[�̨��1���BΜ�@Y�$�q�'f��;�t"���"EAp���	;�0�,�"���5�츐7��8�	mo�ԫ˕=R5�31 x�c���n�4�s6`Z�󥤍4ņ�cn�K.jv�gw�P0��  �L����T���ʗ_}�9�u���k;��Y�%�ZzPF��x�u����$�Ǣ���<cZ��N1������Q�Ù�����^!C��(�/\��1�, zA<�a�>�i�
�u<�`!�?�2@����:l��f�c���EG��WM�F�`?������"�0̎Ev@ZKv���>og��ϗ��6|k �WO!-����YF�*yM�P@���`7��'K`�4��O=H� B Fg��L���g�Y��7���38�g�S��E���k�񊵊muGsJq�qn�tlԃ�ˆCt���3Y$m�"Đ�	��b�M�L�|��u�d��T�\�uE�0��>���S���H��,��X�+�����B���Z��KvT[K<5�=�X�-6e�r�P $�B �Xi.�۝������_9>]�� �]������	{!�b���IkL�`πX�@4tm�1e��,7;Ԥq��e�����	H���n�Vl R�+��/�����9���x�f�8�����]R�k�bS����~W9n=%���EOKx�>c�8�q �'����L�|z���30�ˌ+���1�L4�哶|���m��i�1�4ـ9��]�L8��C�K��p'��Io�	���?��tݨ��R�fC޽8���Am I�h�Qf癘*���	n��Tl����
 � �I��0�o���4V�)� KnMe�i�����F?q����$��V}��׻<�}�ی.�+nT���K۹A �  " ,h �P"�5@H�4 LF!�����AH�-��h�����Ǌt>��F��c��*çB�d�؊��1Q�:����qө��ǅ����9�f�|�Oi��[�s��+��*^��t��1���Vxzf$řp\k�:�|��;�\��U��2C���f1>Dy�"k��������1�f=e8�0�� �r�{�F�.�n4�Jz/��;Q�%���2�TF*
gλg/*I.s�D @����*E$ �l�*@  Y@��R� ��p)u-DUS��p�o�2�iYE��j������
m��6�+���፥����ڱ&v�@J<�M�[^3e-"4�q]�f1�j�#%5�(ɥY�iRJ�8�͉��G9f�E�..�����]��۶A�ҝ��[ˉN5]�$e���#�K�eDK��)4m5�QA�9&um��6q�H�(�J�g��ne�ЁGpƦƶ�����&���R��^$���\�%.:mI3K��0PTRE�<������D��8W��@�~7��l���� ��7w$� �PUx�X�1��J��WLh���,�L�y�b�N�F�Y�1U����,;3uc"��X�l�TS)E�0�#���� 5���Ґ4�c� [b��\�H`��Gs�D��|k�@O��������p��W sA�T��U��V���\.��,�����.�����	!	و}ɸ�f���(k��e[��A0�^!!���i���N�b����O��"��8bN�*V]&�5��#'���<~y����}��U�'IMGH�d�� d�qe��s��*<��O<Ϭ��G��σ�e�-�`=݊u�52a�h����}����#-�&��ڗx4 ��R[�o=ˑ�1o1�!1�Z�T��1��a��zyNa�`�>w��>4%�Ŋ����Dm]{��k�q Ykw��wdO
�UU	���w���@p�%"-��:���>1������E��o�:XA�M�op&�8i���@��ѽ��hZY����`Z"ƌ03�ܻ�9�zyw~�w��3����_%wʠ�j��
�],�T�Xgl��\َ���fj\-���d5#��rB�+�Ť�v����_<錳1����L%eV�԰T��`��'�u��M��d�@�e�L�~p'�-@��\�����B������孒0����4`c32 �:�"b-e�K\���7>{���Οg�'�0�/�����W��DX��P��t_�L<��[��g�ƃK_��%�������{�jj��VmlTD^כ<����sw�����V-]C�^[o�&���"��,sl�d�C���'`il��e_<����Ɠ'ܳ����pZ�XPj�����;����uܥ�voQ0����%X�\;�ލ����V�(��}��ǁ��y�a���a��M�z�s�2JS"Y����	�5ז��}�}s�g�ϟb_[SF�["n���L=1���om�;4�Kz�T�����o���H" �����ff��g_z�>u|9��=��]���s~�
���X�ՕY\�q�2P]E9H,˶���0��9-�A��)*Ie��m��Ap��J�[*�&���mi3e�ew�O+�>W�uuE�0�Cd$4��]zU��M���ߝ��[�À+�U��cV�Fn�qf��s��pF%mÑܠ���~_B���]�o�Ϭ%�s��|��s��A�}0{��Z�㋶���0۳�À������q�k`e�L��2]8���<D�� ��LL���@�����}a�=l<���V-��z�z=��J#q����,���=<�FХ����u�W��ӻ��8�G�nʺT���Z���e�̆$Y6���"���o�o=HM�<��E,0}aG�Sמ$O��7�2j��!Ǽk<P�)�)�R1�d�,/5�br�VS<yb>W�3�!�|�(�׬�dE<��;��ݥ���"��ǓN��w��t�
e��5Ԙ �Ȣ�*X,ND_��S����j��b�W��[oX�G�y��&RRDi�d�Lɦ��SL�IM��Y�)S,ԥ�1T)a�$cE��$	Īi�`E�XČ ��y���e4��ʚRi&l�J2�ͼfi,Sy癱i�L�h�l�0���ȵ�P�̃�5�M�hZ���σ�M�����L�<A��"C��$ΔC���́��0�U���<{��/j���h'�?*��Th��EӠ��t���Y'6%}����4���� =�A��}�1�'*:)�x(��Q�sI��~{䞡;�^����P^���	�������[�n)���C0����<0��^��xh�x1 ;�l��d�n��}M�����������:�,kF��ܥF��&0M��u��s�d�.7f��SFl-"#o)�`�3�j�^ExĨĮa�C�à*�v6�$�޹a����CV�՜�&�
����a�@X� 0�J�X��}1��:31]�\���B*Vf7-��z�9�Nx�4�c���>D��r(��;��W��d��G��Q _	��@� ְ��"ŀ�~�`������Z����*�vY9���\+\-U�
�q;�o+l�Tx�[Ϲ�4����ǉ�}ݐ��7��kȼܷ��dW�=L�����Ŷa�f &��p9�7��~}��7�9���8]����q�dr*��rw�����\�[���P����6����50�:� ø��1q������wc�E: ʧ�x�����^��*��f͂7e��
�Dho5�O�����5n�"�G�;Һ�y�\	�xT�����i�� W���섺�0��E�ˋ]	�nN!�2a���3>|���^.c�d<�3!D�@����M��ܶ$����#�K,�u�h%�FwZ:إ���@��S]�c��2������Iq����0	x���$�y�<����iԧ�m�� ��<;������t[�U|� �|�2oos�5�����Q�-�33,!Bxxvh1ʍ�Z\��~z�w��|��kX��E/J��kán����NT�vl0�-��E0�#v�Ző͍������ O�'{���ZDxN���
I�ࠞ0��@��Ы�Xa^���w��"��ܼ���s�n��{��7�` ſ>3us����j��6��;k��Xd<���F�.��ux���ڈ�:}��׌/Z��i<i��ʃz�n������%u���m��^�j���K�T�iȷ������O�_Rn���T�(-2E�����6I��5���vn���z���޷���s
o8aY�1�}1�k��<������4X�� \�ǜ�y+  _��k�UT(}I� G�׬6R�Ah�lU��_`�~%� g|7	���ǒ��=�!ʞq8�%��\�t��ʿ��� X�+*���)A/mT��r�@��ae��� �R!���bdڊlX,�A�Zb�B �"B"
"B @h�-Eh��N1�L��EQr��c""�6��
�� �x"�a=��  ȡ���V4�5Qm ļ)D�@KDD��Pm@�B�"�rҁj(BH
^7���¤h��n,hY-�X�����m����f�tbª.ZP�-�\��$�IK����BK��%B"(����"����) Hȁ�V��z����K�iP��mmq�eջ�˛���R��i:�)����?���'��rB��C���x����KQ��1��b؄��ւǗ�[rB��V����f�.�N=�$!$�(�z��\�������p�$�!�?K���&��s�ZTP��A��I�d9�(=`@?O�!������	�  G�r2"�~#D ���*Y؁��m�9&��?�jw����y�@z�0v� ����ȅ��RୃJD�n�S7���{��P�Tݼ�5��� e�x ���d�	>�I$�u���Y1��{H_��9��C.���� .�i�,����A0�/\�.V��ȩxFD�Ry-�5>;���������� �qLR����7�;��L��c������v�&�e�KS�������
�b/AxV�����$w�oP mW�E��
 -���0N*�o��\0Ȓ
�!�(����FZR��H"� "U�R�6$����EkQb�X���F�a�1` A��@�E�B#( @dA	 A" � �	$AdVEd@�*
E��b�X��X�����"$U�œd�K,�Y6f��Jb��"Ȭ ��`�� @.@UP��� �"(�Ci�Q`"FD"�\-���±ԣ4����{��V�ݶ�P�.�?:xz�FH�u��/A3 G�t �Yc�f}9���p�ǥ���r�����R�%XMS�J����^���s;z��Oô�d�f���Q�7V��y)ۦ�H���ʞ=��}=�p�������z~]l�Љ�yO��lf�JsK���$��E�4XѢƍQ4X�bƋ4�h�cFƍMѢƋ,XѢ4h�b�E�,F͕*664XѢ4TX�,�-Zh�,�,ѳe��4F�4Y4h��FѣE��4Xѣ��fh��E�%4h��ƍ�lh�#F���cF���#EIcL���cF�M-4�4XѢƋ�f͍)XѢƚh�,TZ4�f�Di,�4�4XѢ4h�4YK,h�#F�,�,Y,�"4�j,i,i�,h�F�2��cF�F��bƍ�,h؍F�,Xѱ�E,j4X��Ţ�h�cE�,h�#F�*-,h�4Y66M&�4cF��E�K6#F�kK)�E�F�$�&�,h�cI�,�QcE�,���R�lXѱcE�2h���cF�I4h��Q�4YK&h�cFƋ,K4h�b�Ƌ,��E����64F�,X�X�XѴh�d�dѢƍ���h�h�4h��E3I�Ƌ,li4F�2ƍ�,i,I�E�fŢɣD�4Y,li,Y4X���ɢƍ4h�F�ƒƍ4L��l��h�M�4F��ƒŒ�dѣ6,h���I�ّLѢƒ�cbƋ�E�4YM�#L�Y�*4X��F�,X�X�Q�I4X�cF�#F�M�64�#cIcE�,�$Ѣɱ�h�Q�I%�%�4i,X�4X�d��d�b#EIb�cF�&��cḇ��Ƌ�,Xѱ��ɣIM4�,�,h�4͍4h��؍&�K6,h�M4X�d�d�4k&�cE�Ƌ�IQbɴh���$�Xٚ,X�,h�$X�Xѱ��ƓF�,h�S4X�b�,�*4���I��!������Ɉ�IQ�(��J02ABA�dI�d����
 E��b'!�����6;�33��X�C�}r�RiY�����KQ�g�c3��dbz��.N[������^5�M�u�H�+��2w����qb��,;>�2C��R{��/�L�)�y�|����!���_!ET��Lbb ��R�ܞ
Cܞqd�c�c3��z�1z�R��v�ĆϜ|��x���� ����&]t*�K�1g�<݁���h��zrY*�^e�Bxq�D:��C�E��li�&�`���K��L�=�u�  ��C4���JP~���C�b�$�.'� ��)ָ'q@�����Id�J�
�宲A.�
��a���Gww��"OV����X�%��Ղ֨T����X ����r�	��EGD�`�)0�.R�*�^i�� fP��.���2�-B�0��.:.Рꤌ(aj��@JQ[��yTA:fk��� ��_�p��(���ڞ�3W�Ag��+�Lw��DU>�s̱M`/'���~b~�����p�/7��[����tR���==�n��"y��'rz�<��#�#���{"`���B���f�bs��d/؜ƅP6/t�;�A�THH]jఉ/2��R#1����(�*{ۂ�(bi�\KF����� ��0^���`h�i 􁚙�&��܃�m`�v��za��iD!QU!0�� ���&�$���L���D�3O@9�.����\/~&��VAb,(�pNFZ��f.�,�=jm���q8��I$�Q�9�0M?�������/\���Z�K@;@��0�TI��I%��6Ɂ49�ȭ"]�'$�!+ږ���dqX&!���3������l�%��GU��SF%%�֪����F�sM��2�60A�[��w;Q�~��F�sg儋��=�G���M{{�UA���Q@=��|�B����J�%�|w�.���pw
��МǠ�ax����ú��K�)�m�23�5�M�"eZD��>1?��S�#�G/E�����g���/iЮY8	=�H��`A�����w$S�	��E�